magic
tech sky130A
timestamp 1654591597
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4365 -480 4421 240
rect 4963 -480 5019 240
rect 5561 -480 5617 240
rect 6159 -480 6215 240
rect 6757 -480 6813 240
rect 7355 -480 7411 240
rect 7953 -480 8009 240
rect 8505 -480 8561 240
rect 9103 -480 9159 240
rect 9701 -480 9757 240
rect 10299 -480 10355 240
rect 10897 -480 10953 240
rect 11495 -480 11551 240
rect 12093 -480 12149 240
rect 12645 -480 12701 240
rect 13243 -480 13299 240
rect 13841 -480 13897 240
rect 14439 -480 14495 240
rect 15037 -480 15093 240
rect 15635 -480 15691 240
rect 16187 -480 16243 240
rect 16785 -480 16841 240
rect 17383 -480 17439 240
rect 17981 -480 18037 240
rect 18579 -480 18635 240
rect 19177 -480 19233 240
rect 19775 -480 19831 240
rect 20327 -480 20383 240
rect 20925 -480 20981 240
rect 21523 -480 21579 240
rect 22121 -480 22177 240
rect 22719 -480 22775 240
rect 23317 -480 23373 240
rect 23915 -480 23971 240
rect 24467 -480 24523 240
rect 25065 -480 25121 240
rect 25663 -480 25719 240
rect 26261 -480 26317 240
rect 26859 -480 26915 240
rect 27457 -480 27513 240
rect 28009 -480 28065 240
rect 28607 -480 28663 240
rect 29205 -480 29261 240
rect 29803 -480 29859 240
rect 30401 -480 30457 240
rect 30999 -480 31055 240
rect 31597 -480 31653 240
rect 32149 -480 32205 240
rect 32747 -480 32803 240
rect 33345 -480 33401 240
rect 33943 -480 33999 240
rect 34541 -480 34597 240
rect 35139 -480 35195 240
rect 35737 -480 35793 240
rect 36289 -480 36345 240
rect 36887 -480 36943 240
rect 37485 -480 37541 240
rect 38083 -480 38139 240
rect 38681 -480 38737 240
rect 39279 -480 39335 240
rect 39831 -480 39887 240
rect 40429 -480 40485 240
rect 41027 -480 41083 240
rect 41625 -480 41681 240
rect 42223 -480 42279 240
rect 42821 -480 42877 240
rect 43419 -480 43475 240
rect 43971 -480 44027 240
rect 44569 -480 44625 240
rect 45167 -480 45223 240
rect 45765 -480 45821 240
rect 46363 -480 46419 240
rect 46961 -480 47017 240
rect 47559 -480 47615 240
rect 48111 -480 48167 240
rect 48709 -480 48765 240
rect 49307 -480 49363 240
rect 49905 -480 49961 240
rect 50503 -480 50559 240
rect 51101 -480 51157 240
rect 51653 -480 51709 240
rect 52251 -480 52307 240
rect 52849 -480 52905 240
rect 53447 -480 53503 240
rect 54045 -480 54101 240
rect 54643 -480 54699 240
rect 55241 -480 55297 240
rect 55793 -480 55849 240
rect 56391 -480 56447 240
rect 56989 -480 57045 240
rect 57587 -480 57643 240
rect 58185 -480 58241 240
rect 58783 -480 58839 240
rect 59381 -480 59437 240
rect 59933 -480 59989 240
rect 60531 -480 60587 240
rect 61129 -480 61185 240
rect 61727 -480 61783 240
rect 62325 -480 62381 240
rect 62923 -480 62979 240
rect 63475 -480 63531 240
rect 64073 -480 64129 240
rect 64671 -480 64727 240
rect 65269 -480 65325 240
rect 65867 -480 65923 240
rect 66465 -480 66521 240
rect 67063 -480 67119 240
rect 67615 -480 67671 240
rect 68213 -480 68269 240
rect 68811 -480 68867 240
rect 69409 -480 69465 240
rect 70007 -480 70063 240
rect 70605 -480 70661 240
rect 71203 -480 71259 240
rect 71755 -480 71811 240
rect 72353 -480 72409 240
rect 72951 -480 73007 240
rect 73549 -480 73605 240
rect 74147 -480 74203 240
rect 74745 -480 74801 240
rect 75297 -480 75353 240
rect 75895 -480 75951 240
rect 76493 -480 76549 240
rect 77091 -480 77147 240
rect 77689 -480 77745 240
rect 78287 -480 78343 240
rect 78885 -480 78941 240
rect 79437 -480 79493 240
rect 80035 -480 80091 240
rect 80633 -480 80689 240
rect 81231 -480 81287 240
rect 81829 -480 81885 240
rect 82427 -480 82483 240
rect 83025 -480 83081 240
rect 83577 -480 83633 240
rect 84175 -480 84231 240
rect 84773 -480 84829 240
rect 85371 -480 85427 240
rect 85969 -480 86025 240
rect 86567 -480 86623 240
rect 87119 -480 87175 240
rect 87717 -480 87773 240
rect 88315 -480 88371 240
rect 88913 -480 88969 240
rect 89511 -480 89567 240
rect 90109 -480 90165 240
rect 90707 -480 90763 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92455 -480 92511 240
rect 93053 -480 93109 240
rect 93651 -480 93707 240
rect 94249 -480 94305 240
rect 94847 -480 94903 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98941 -480 98997 240
rect 99539 -480 99595 240
rect 100137 -480 100193 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103081 -480 103137 240
rect 103679 -480 103735 240
rect 104277 -480 104333 240
rect 104875 -480 104931 240
rect 105473 -480 105529 240
rect 106071 -480 106127 240
rect 106669 -480 106725 240
rect 107221 -480 107277 240
rect 107819 -480 107875 240
rect 108417 -480 108473 240
rect 109015 -480 109071 240
rect 109613 -480 109669 240
rect 110211 -480 110267 240
rect 110763 -480 110819 240
rect 111361 -480 111417 240
rect 111959 -480 112015 240
rect 112557 -480 112613 240
rect 113155 -480 113211 240
rect 113753 -480 113809 240
rect 114351 -480 114407 240
rect 114903 -480 114959 240
rect 115501 -480 115557 240
rect 116099 -480 116155 240
rect 116697 -480 116753 240
rect 117295 -480 117351 240
rect 117893 -480 117949 240
rect 118491 -480 118547 240
rect 119043 -480 119099 240
rect 119641 -480 119697 240
rect 120239 -480 120295 240
rect 120837 -480 120893 240
rect 121435 -480 121491 240
rect 122033 -480 122089 240
rect 122585 -480 122641 240
rect 123183 -480 123239 240
rect 123781 -480 123837 240
rect 124379 -480 124435 240
rect 124977 -480 125033 240
rect 125575 -480 125631 240
rect 126173 -480 126229 240
rect 126725 -480 126781 240
rect 127323 -480 127379 240
rect 127921 -480 127977 240
rect 128519 -480 128575 240
rect 129117 -480 129173 240
rect 129715 -480 129771 240
rect 130313 -480 130369 240
rect 130865 -480 130921 240
rect 131463 -480 131519 240
rect 132061 -480 132117 240
rect 132659 -480 132715 240
rect 133257 -480 133313 240
rect 133855 -480 133911 240
rect 134407 -480 134463 240
rect 135005 -480 135061 240
rect 135603 -480 135659 240
rect 136201 -480 136257 240
rect 136799 -480 136855 240
rect 137397 -480 137453 240
rect 137995 -480 138051 240
rect 138547 -480 138603 240
rect 139145 -480 139201 240
rect 139743 -480 139799 240
rect 140341 -480 140397 240
rect 140939 -480 140995 240
rect 141537 -480 141593 240
rect 142135 -480 142191 240
rect 142687 -480 142743 240
rect 143285 -480 143341 240
rect 143883 -480 143939 240
rect 144481 -480 144537 240
rect 145079 -480 145135 240
rect 145677 -480 145733 240
rect 146275 -480 146331 240
rect 146827 -480 146883 240
rect 147425 -480 147481 240
rect 148023 -480 148079 240
rect 148621 -480 148677 240
rect 149219 -480 149275 240
rect 149817 -480 149873 240
rect 150369 -480 150425 240
rect 150967 -480 151023 240
rect 151565 -480 151621 240
rect 152163 -480 152219 240
rect 152761 -480 152817 240
rect 153359 -480 153415 240
rect 153957 -480 154013 240
rect 154509 -480 154565 240
rect 155107 -480 155163 240
rect 155705 -480 155761 240
rect 156303 -480 156359 240
rect 156901 -480 156957 240
rect 157499 -480 157555 240
rect 158097 -480 158153 240
rect 158649 -480 158705 240
rect 159247 -480 159303 240
rect 159845 -480 159901 240
rect 160443 -480 160499 240
rect 161041 -480 161097 240
rect 161639 -480 161695 240
rect 162191 -480 162247 240
rect 162789 -480 162845 240
rect 163387 -480 163443 240
rect 163985 -480 164041 240
rect 164583 -480 164639 240
rect 165181 -480 165237 240
rect 165779 -480 165835 240
rect 166331 -480 166387 240
rect 166929 -480 166985 240
rect 167527 -480 167583 240
rect 168125 -480 168181 240
rect 168723 -480 168779 240
rect 169321 -480 169377 240
rect 169919 -480 169975 240
rect 170471 -480 170527 240
rect 171069 -480 171125 240
rect 171667 -480 171723 240
rect 172265 -480 172321 240
rect 172863 -480 172919 240
rect 173461 -480 173517 240
rect 174013 -480 174069 240
rect 174611 -480 174667 240
rect 175209 -480 175265 240
rect 175807 -480 175863 240
rect 176405 -480 176461 240
rect 177003 -480 177059 240
rect 177601 -480 177657 240
rect 178153 -480 178209 240
rect 178751 -480 178807 240
rect 179349 -480 179405 240
rect 179947 -480 180003 240
rect 180545 -480 180601 240
rect 181143 -480 181199 240
rect 181741 -480 181797 240
rect 182293 -480 182349 240
rect 182891 -480 182947 240
rect 183489 -480 183545 240
rect 184087 -480 184143 240
rect 184685 -480 184741 240
rect 185283 -480 185339 240
rect 185835 -480 185891 240
rect 186433 -480 186489 240
rect 187031 -480 187087 240
rect 187629 -480 187685 240
rect 188227 -480 188283 240
rect 188825 -480 188881 240
rect 189423 -480 189479 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192367 -480 192423 240
rect 192965 -480 193021 240
rect 193563 -480 193619 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197657 -480 197713 240
rect 198255 -480 198311 240
rect 198853 -480 198909 240
rect 199451 -480 199507 240
rect 200049 -480 200105 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201797 -480 201853 240
rect 202395 -480 202451 240
rect 202993 -480 203049 240
rect 203591 -480 203647 240
rect 204189 -480 204245 240
rect 204787 -480 204843 240
rect 205385 -480 205441 240
rect 205937 -480 205993 240
rect 206535 -480 206591 240
rect 207133 -480 207189 240
rect 207731 -480 207787 240
rect 208329 -480 208385 240
rect 208927 -480 208983 240
rect 209479 -480 209535 240
rect 210077 -480 210133 240
rect 210675 -480 210731 240
rect 211273 -480 211329 240
rect 211871 -480 211927 240
rect 212469 -480 212525 240
rect 213067 -480 213123 240
rect 213619 -480 213675 240
rect 214217 -480 214273 240
rect 214815 -480 214871 240
rect 215413 -480 215469 240
rect 216011 -480 216067 240
rect 216609 -480 216665 240
rect 217207 -480 217263 240
rect 217759 -480 217815 240
rect 218357 -480 218413 240
rect 218955 -480 219011 240
rect 219553 -480 219609 240
rect 220151 -480 220207 240
rect 220749 -480 220805 240
rect 221301 -480 221357 240
rect 221899 -480 221955 240
rect 222497 -480 222553 240
rect 223095 -480 223151 240
rect 223693 -480 223749 240
rect 224291 -480 224347 240
rect 224889 -480 224945 240
rect 225441 -480 225497 240
rect 226039 -480 226095 240
rect 226637 -480 226693 240
rect 227235 -480 227291 240
rect 227833 -480 227889 240
rect 228431 -480 228487 240
rect 229029 -480 229085 240
rect 229581 -480 229637 240
rect 230179 -480 230235 240
rect 230777 -480 230833 240
rect 231375 -480 231431 240
rect 231973 -480 232029 240
rect 232571 -480 232627 240
rect 233123 -480 233179 240
rect 233721 -480 233777 240
rect 234319 -480 234375 240
rect 234917 -480 234973 240
rect 235515 -480 235571 240
rect 236113 -480 236169 240
rect 236711 -480 236767 240
rect 237263 -480 237319 240
rect 237861 -480 237917 240
rect 238459 -480 238515 240
rect 239057 -480 239113 240
rect 239655 -480 239711 240
rect 240253 -480 240309 240
rect 240851 -480 240907 240
rect 241403 -480 241459 240
rect 242001 -480 242057 240
rect 242599 -480 242655 240
rect 243197 -480 243253 240
rect 243795 -480 243851 240
rect 244393 -480 244449 240
rect 244945 -480 245001 240
rect 245543 -480 245599 240
rect 246141 -480 246197 240
rect 246739 -480 246795 240
rect 247337 -480 247393 240
rect 247935 -480 247991 240
rect 248533 -480 248589 240
rect 249085 -480 249141 240
rect 249683 -480 249739 240
rect 250281 -480 250337 240
rect 250879 -480 250935 240
rect 251477 -480 251533 240
rect 252075 -480 252131 240
rect 252673 -480 252729 240
rect 253225 -480 253281 240
rect 253823 -480 253879 240
rect 254421 -480 254477 240
rect 255019 -480 255075 240
rect 255617 -480 255673 240
rect 256215 -480 256271 240
rect 256767 -480 256823 240
rect 257365 -480 257421 240
rect 257963 -480 258019 240
rect 258561 -480 258617 240
rect 259159 -480 259215 240
rect 259757 -480 259813 240
rect 260355 -480 260411 240
rect 260907 -480 260963 240
rect 261505 -480 261561 240
rect 262103 -480 262159 240
rect 262701 -480 262757 240
rect 263299 -480 263355 240
rect 263897 -480 263953 240
rect 264495 -480 264551 240
rect 265047 -480 265103 240
rect 265645 -480 265701 240
rect 266243 -480 266299 240
rect 266841 -480 266897 240
rect 267439 -480 267495 240
rect 268037 -480 268093 240
rect 268589 -480 268645 240
rect 269187 -480 269243 240
rect 269785 -480 269841 240
rect 270383 -480 270439 240
rect 270981 -480 271037 240
rect 271579 -480 271635 240
rect 272177 -480 272233 240
rect 272729 -480 272785 240
rect 273327 -480 273383 240
rect 273925 -480 273981 240
rect 274523 -480 274579 240
rect 275121 -480 275177 240
rect 275719 -480 275775 240
rect 276317 -480 276373 240
rect 276869 -480 276925 240
rect 277467 -480 277523 240
rect 278065 -480 278121 240
rect 278663 -480 278719 240
rect 279261 -480 279317 240
rect 279859 -480 279915 240
rect 280411 -480 280467 240
rect 281009 -480 281065 240
rect 281607 -480 281663 240
rect 282205 -480 282261 240
rect 282803 -480 282859 240
rect 283401 -480 283457 240
rect 283999 -480 284055 240
rect 284551 -480 284607 240
rect 285149 -480 285205 240
rect 285747 -480 285803 240
rect 286345 -480 286401 240
rect 286943 -480 286999 240
rect 287541 -480 287597 240
rect 288139 -480 288195 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect -480 348610 240 348730
rect 291760 348542 292480 348662
rect -480 342082 240 342202
rect 291760 341878 292480 341998
rect -480 335554 240 335674
rect 291760 335282 292480 335402
rect -480 329026 240 329146
rect 291760 328618 292480 328738
rect -480 322498 240 322618
rect 291760 321954 292480 322074
rect -480 315970 240 316090
rect 291760 315358 292480 315478
rect -480 309510 240 309630
rect 291760 308694 292480 308814
rect -480 302982 240 303102
rect 291760 302030 292480 302150
rect -480 296454 240 296574
rect 291760 295434 292480 295554
rect -480 289926 240 290046
rect 291760 288770 292480 288890
rect -480 283398 240 283518
rect 291760 282106 292480 282226
rect -480 276870 240 276990
rect 291760 275510 292480 275630
rect -480 270342 240 270462
rect 291760 268846 292480 268966
rect -480 263882 240 264002
rect 291760 262182 292480 262302
rect -480 257354 240 257474
rect 291760 255586 292480 255706
rect -480 250826 240 250946
rect 291760 248922 292480 249042
rect -480 244298 240 244418
rect 291760 242258 292480 242378
rect -480 237770 240 237890
rect 291760 235662 292480 235782
rect -480 231242 240 231362
rect 291760 228998 292480 229118
rect -480 224714 240 224834
rect 291760 222334 292480 222454
rect -480 218254 240 218374
rect 291760 215738 292480 215858
rect -480 211726 240 211846
rect 291760 209074 292480 209194
rect -480 205198 240 205318
rect 291760 202410 292480 202530
rect -480 198670 240 198790
rect 291760 195814 292480 195934
rect -480 192142 240 192262
rect 291760 189150 292480 189270
rect -480 185614 240 185734
rect 291760 182486 292480 182606
rect -480 179154 240 179274
rect 291760 175890 292480 176010
rect -480 172626 240 172746
rect 291760 169226 292480 169346
rect -480 166098 240 166218
rect 291760 162562 292480 162682
rect -480 159570 240 159690
rect 291760 155966 292480 156086
rect -480 153042 240 153162
rect 291760 149302 292480 149422
rect -480 146514 240 146634
rect 291760 142638 292480 142758
rect -480 139986 240 140106
rect 291760 136042 292480 136162
rect -480 133526 240 133646
rect 291760 129378 292480 129498
rect -480 126998 240 127118
rect 291760 122714 292480 122834
rect -480 120470 240 120590
rect 291760 116118 292480 116238
rect -480 113942 240 114062
rect 291760 109454 292480 109574
rect -480 107414 240 107534
rect 291760 102790 292480 102910
rect -480 100886 240 101006
rect 291760 96194 292480 96314
rect -480 94358 240 94478
rect 291760 89530 292480 89650
rect -480 87898 240 88018
rect 291760 82866 292480 82986
rect -480 81370 240 81490
rect 291760 76270 292480 76390
rect -480 74842 240 74962
rect 291760 69606 292480 69726
rect -480 68314 240 68434
rect 291760 62942 292480 63062
rect -480 61786 240 61906
rect 291760 56346 292480 56466
rect -480 55258 240 55378
rect 291760 49682 292480 49802
rect -480 48730 240 48850
rect 291760 43018 292480 43138
rect -480 42270 240 42390
rect 291760 36422 292480 36542
rect -480 35742 240 35862
rect 291760 29758 292480 29878
rect -480 29214 240 29334
rect 291760 23094 292480 23214
rect -480 22686 240 22806
rect 291760 16498 292480 16618
rect -480 16158 240 16278
rect 291760 9834 292480 9954
rect -480 9630 240 9750
rect -480 3170 240 3290
rect 291760 3238 292480 3358
<< metal4 >>
rect -4363 355779 -4053 355795
rect -4363 355501 -4347 355779
rect -4069 355501 -4053 355779
rect -4363 340307 -4053 355501
rect -4363 340029 -4347 340307
rect -4069 340029 -4053 340307
rect -4363 322307 -4053 340029
rect -4363 322029 -4347 322307
rect -4069 322029 -4053 322307
rect -4363 304307 -4053 322029
rect -4363 304029 -4347 304307
rect -4069 304029 -4053 304307
rect -4363 286307 -4053 304029
rect -4363 286029 -4347 286307
rect -4069 286029 -4053 286307
rect -4363 268307 -4053 286029
rect -4363 268029 -4347 268307
rect -4069 268029 -4053 268307
rect -4363 250307 -4053 268029
rect -4363 250029 -4347 250307
rect -4069 250029 -4053 250307
rect -4363 232307 -4053 250029
rect -4363 232029 -4347 232307
rect -4069 232029 -4053 232307
rect -4363 214307 -4053 232029
rect -4363 214029 -4347 214307
rect -4069 214029 -4053 214307
rect -4363 196307 -4053 214029
rect -4363 196029 -4347 196307
rect -4069 196029 -4053 196307
rect -4363 178307 -4053 196029
rect -4363 178029 -4347 178307
rect -4069 178029 -4053 178307
rect -4363 160307 -4053 178029
rect -4363 160029 -4347 160307
rect -4069 160029 -4053 160307
rect -4363 142307 -4053 160029
rect -4363 142029 -4347 142307
rect -4069 142029 -4053 142307
rect -4363 124307 -4053 142029
rect -4363 124029 -4347 124307
rect -4069 124029 -4053 124307
rect -4363 106307 -4053 124029
rect -4363 106029 -4347 106307
rect -4069 106029 -4053 106307
rect -4363 88307 -4053 106029
rect -4363 88029 -4347 88307
rect -4069 88029 -4053 88307
rect -4363 70307 -4053 88029
rect -4363 70029 -4347 70307
rect -4069 70029 -4053 70307
rect -4363 52307 -4053 70029
rect -4363 52029 -4347 52307
rect -4069 52029 -4053 52307
rect -4363 34307 -4053 52029
rect -4363 34029 -4347 34307
rect -4069 34029 -4053 34307
rect -4363 16307 -4053 34029
rect -4363 16029 -4347 16307
rect -4069 16029 -4053 16307
rect -4363 -3533 -4053 16029
rect -3883 355299 -3573 355315
rect -3883 355021 -3867 355299
rect -3589 355021 -3573 355299
rect -3883 349307 -3573 355021
rect 6477 355299 6787 355795
rect 6477 355021 6493 355299
rect 6771 355021 6787 355299
rect -3883 349029 -3867 349307
rect -3589 349029 -3573 349307
rect -3883 331307 -3573 349029
rect -3883 331029 -3867 331307
rect -3589 331029 -3573 331307
rect -3883 313307 -3573 331029
rect -3883 313029 -3867 313307
rect -3589 313029 -3573 313307
rect -3883 295307 -3573 313029
rect -3883 295029 -3867 295307
rect -3589 295029 -3573 295307
rect -3883 277307 -3573 295029
rect -3883 277029 -3867 277307
rect -3589 277029 -3573 277307
rect -3883 259307 -3573 277029
rect -3883 259029 -3867 259307
rect -3589 259029 -3573 259307
rect -3883 241307 -3573 259029
rect -3883 241029 -3867 241307
rect -3589 241029 -3573 241307
rect -3883 223307 -3573 241029
rect -3883 223029 -3867 223307
rect -3589 223029 -3573 223307
rect -3883 205307 -3573 223029
rect -3883 205029 -3867 205307
rect -3589 205029 -3573 205307
rect -3883 187307 -3573 205029
rect -3883 187029 -3867 187307
rect -3589 187029 -3573 187307
rect -3883 169307 -3573 187029
rect -3883 169029 -3867 169307
rect -3589 169029 -3573 169307
rect -3883 151307 -3573 169029
rect -3883 151029 -3867 151307
rect -3589 151029 -3573 151307
rect -3883 133307 -3573 151029
rect -3883 133029 -3867 133307
rect -3589 133029 -3573 133307
rect -3883 115307 -3573 133029
rect -3883 115029 -3867 115307
rect -3589 115029 -3573 115307
rect -3883 97307 -3573 115029
rect -3883 97029 -3867 97307
rect -3589 97029 -3573 97307
rect -3883 79307 -3573 97029
rect -3883 79029 -3867 79307
rect -3589 79029 -3573 79307
rect -3883 61307 -3573 79029
rect -3883 61029 -3867 61307
rect -3589 61029 -3573 61307
rect -3883 43307 -3573 61029
rect -3883 43029 -3867 43307
rect -3589 43029 -3573 43307
rect -3883 25307 -3573 43029
rect -3883 25029 -3867 25307
rect -3589 25029 -3573 25307
rect -3883 7307 -3573 25029
rect -3883 7029 -3867 7307
rect -3589 7029 -3573 7307
rect -3883 -3053 -3573 7029
rect -3403 354819 -3093 354835
rect -3403 354541 -3387 354819
rect -3109 354541 -3093 354819
rect -3403 338447 -3093 354541
rect -3403 338169 -3387 338447
rect -3109 338169 -3093 338447
rect -3403 320447 -3093 338169
rect -3403 320169 -3387 320447
rect -3109 320169 -3093 320447
rect -3403 302447 -3093 320169
rect -3403 302169 -3387 302447
rect -3109 302169 -3093 302447
rect -3403 284447 -3093 302169
rect -3403 284169 -3387 284447
rect -3109 284169 -3093 284447
rect -3403 266447 -3093 284169
rect -3403 266169 -3387 266447
rect -3109 266169 -3093 266447
rect -3403 248447 -3093 266169
rect -3403 248169 -3387 248447
rect -3109 248169 -3093 248447
rect -3403 230447 -3093 248169
rect -3403 230169 -3387 230447
rect -3109 230169 -3093 230447
rect -3403 212447 -3093 230169
rect -3403 212169 -3387 212447
rect -3109 212169 -3093 212447
rect -3403 194447 -3093 212169
rect -3403 194169 -3387 194447
rect -3109 194169 -3093 194447
rect -3403 176447 -3093 194169
rect -3403 176169 -3387 176447
rect -3109 176169 -3093 176447
rect -3403 158447 -3093 176169
rect -3403 158169 -3387 158447
rect -3109 158169 -3093 158447
rect -3403 140447 -3093 158169
rect -3403 140169 -3387 140447
rect -3109 140169 -3093 140447
rect -3403 122447 -3093 140169
rect -3403 122169 -3387 122447
rect -3109 122169 -3093 122447
rect -3403 104447 -3093 122169
rect -3403 104169 -3387 104447
rect -3109 104169 -3093 104447
rect -3403 86447 -3093 104169
rect -3403 86169 -3387 86447
rect -3109 86169 -3093 86447
rect -3403 68447 -3093 86169
rect -3403 68169 -3387 68447
rect -3109 68169 -3093 68447
rect -3403 50447 -3093 68169
rect -3403 50169 -3387 50447
rect -3109 50169 -3093 50447
rect -3403 32447 -3093 50169
rect -3403 32169 -3387 32447
rect -3109 32169 -3093 32447
rect -3403 14447 -3093 32169
rect -3403 14169 -3387 14447
rect -3109 14169 -3093 14447
rect -3403 -2573 -3093 14169
rect -2923 354339 -2613 354355
rect -2923 354061 -2907 354339
rect -2629 354061 -2613 354339
rect -2923 347447 -2613 354061
rect 4617 354339 4927 354835
rect 4617 354061 4633 354339
rect 4911 354061 4927 354339
rect -2923 347169 -2907 347447
rect -2629 347169 -2613 347447
rect -2923 329447 -2613 347169
rect -2923 329169 -2907 329447
rect -2629 329169 -2613 329447
rect -2923 311447 -2613 329169
rect -2923 311169 -2907 311447
rect -2629 311169 -2613 311447
rect -2923 293447 -2613 311169
rect -2923 293169 -2907 293447
rect -2629 293169 -2613 293447
rect -2923 275447 -2613 293169
rect -2923 275169 -2907 275447
rect -2629 275169 -2613 275447
rect -2923 257447 -2613 275169
rect -2923 257169 -2907 257447
rect -2629 257169 -2613 257447
rect -2923 239447 -2613 257169
rect -2923 239169 -2907 239447
rect -2629 239169 -2613 239447
rect -2923 221447 -2613 239169
rect -2923 221169 -2907 221447
rect -2629 221169 -2613 221447
rect -2923 203447 -2613 221169
rect -2923 203169 -2907 203447
rect -2629 203169 -2613 203447
rect -2923 185447 -2613 203169
rect -2923 185169 -2907 185447
rect -2629 185169 -2613 185447
rect -2923 167447 -2613 185169
rect -2923 167169 -2907 167447
rect -2629 167169 -2613 167447
rect -2923 149447 -2613 167169
rect -2923 149169 -2907 149447
rect -2629 149169 -2613 149447
rect -2923 131447 -2613 149169
rect -2923 131169 -2907 131447
rect -2629 131169 -2613 131447
rect -2923 113447 -2613 131169
rect -2923 113169 -2907 113447
rect -2629 113169 -2613 113447
rect -2923 95447 -2613 113169
rect -2923 95169 -2907 95447
rect -2629 95169 -2613 95447
rect -2923 77447 -2613 95169
rect -2923 77169 -2907 77447
rect -2629 77169 -2613 77447
rect -2923 59447 -2613 77169
rect -2923 59169 -2907 59447
rect -2629 59169 -2613 59447
rect -2923 41447 -2613 59169
rect -2923 41169 -2907 41447
rect -2629 41169 -2613 41447
rect -2923 23447 -2613 41169
rect -2923 23169 -2907 23447
rect -2629 23169 -2613 23447
rect -2923 5447 -2613 23169
rect -2923 5169 -2907 5447
rect -2629 5169 -2613 5447
rect -2923 -2093 -2613 5169
rect -2443 353859 -2133 353875
rect -2443 353581 -2427 353859
rect -2149 353581 -2133 353859
rect -2443 336587 -2133 353581
rect -2443 336309 -2427 336587
rect -2149 336309 -2133 336587
rect -2443 318587 -2133 336309
rect -2443 318309 -2427 318587
rect -2149 318309 -2133 318587
rect -2443 300587 -2133 318309
rect -2443 300309 -2427 300587
rect -2149 300309 -2133 300587
rect -2443 282587 -2133 300309
rect -2443 282309 -2427 282587
rect -2149 282309 -2133 282587
rect -2443 264587 -2133 282309
rect -2443 264309 -2427 264587
rect -2149 264309 -2133 264587
rect -2443 246587 -2133 264309
rect -2443 246309 -2427 246587
rect -2149 246309 -2133 246587
rect -2443 228587 -2133 246309
rect -2443 228309 -2427 228587
rect -2149 228309 -2133 228587
rect -2443 210587 -2133 228309
rect -2443 210309 -2427 210587
rect -2149 210309 -2133 210587
rect -2443 192587 -2133 210309
rect -2443 192309 -2427 192587
rect -2149 192309 -2133 192587
rect -2443 174587 -2133 192309
rect -2443 174309 -2427 174587
rect -2149 174309 -2133 174587
rect -2443 156587 -2133 174309
rect -2443 156309 -2427 156587
rect -2149 156309 -2133 156587
rect -2443 138587 -2133 156309
rect -2443 138309 -2427 138587
rect -2149 138309 -2133 138587
rect -2443 120587 -2133 138309
rect -2443 120309 -2427 120587
rect -2149 120309 -2133 120587
rect -2443 102587 -2133 120309
rect -2443 102309 -2427 102587
rect -2149 102309 -2133 102587
rect -2443 84587 -2133 102309
rect -2443 84309 -2427 84587
rect -2149 84309 -2133 84587
rect -2443 66587 -2133 84309
rect -2443 66309 -2427 66587
rect -2149 66309 -2133 66587
rect -2443 48587 -2133 66309
rect -2443 48309 -2427 48587
rect -2149 48309 -2133 48587
rect -2443 30587 -2133 48309
rect -2443 30309 -2427 30587
rect -2149 30309 -2133 30587
rect -2443 12587 -2133 30309
rect -2443 12309 -2427 12587
rect -2149 12309 -2133 12587
rect -2443 -1613 -2133 12309
rect -1963 353379 -1653 353395
rect -1963 353101 -1947 353379
rect -1669 353101 -1653 353379
rect -1963 345587 -1653 353101
rect 2757 353379 3067 353875
rect 2757 353101 2773 353379
rect 3051 353101 3067 353379
rect -1963 345309 -1947 345587
rect -1669 345309 -1653 345587
rect -1963 327587 -1653 345309
rect -1963 327309 -1947 327587
rect -1669 327309 -1653 327587
rect -1963 309587 -1653 327309
rect -1963 309309 -1947 309587
rect -1669 309309 -1653 309587
rect -1963 291587 -1653 309309
rect -1963 291309 -1947 291587
rect -1669 291309 -1653 291587
rect -1963 273587 -1653 291309
rect -1963 273309 -1947 273587
rect -1669 273309 -1653 273587
rect -1963 255587 -1653 273309
rect -1963 255309 -1947 255587
rect -1669 255309 -1653 255587
rect -1963 237587 -1653 255309
rect -1963 237309 -1947 237587
rect -1669 237309 -1653 237587
rect -1963 219587 -1653 237309
rect -1963 219309 -1947 219587
rect -1669 219309 -1653 219587
rect -1963 201587 -1653 219309
rect -1963 201309 -1947 201587
rect -1669 201309 -1653 201587
rect -1963 183587 -1653 201309
rect -1963 183309 -1947 183587
rect -1669 183309 -1653 183587
rect -1963 165587 -1653 183309
rect -1963 165309 -1947 165587
rect -1669 165309 -1653 165587
rect -1963 147587 -1653 165309
rect -1963 147309 -1947 147587
rect -1669 147309 -1653 147587
rect -1963 129587 -1653 147309
rect -1963 129309 -1947 129587
rect -1669 129309 -1653 129587
rect -1963 111587 -1653 129309
rect -1963 111309 -1947 111587
rect -1669 111309 -1653 111587
rect -1963 93587 -1653 111309
rect -1963 93309 -1947 93587
rect -1669 93309 -1653 93587
rect -1963 75587 -1653 93309
rect -1963 75309 -1947 75587
rect -1669 75309 -1653 75587
rect -1963 57587 -1653 75309
rect -1963 57309 -1947 57587
rect -1669 57309 -1653 57587
rect -1963 39587 -1653 57309
rect -1963 39309 -1947 39587
rect -1669 39309 -1653 39587
rect -1963 21587 -1653 39309
rect -1963 21309 -1947 21587
rect -1669 21309 -1653 21587
rect -1963 3587 -1653 21309
rect -1963 3309 -1947 3587
rect -1669 3309 -1653 3587
rect -1963 -1133 -1653 3309
rect -1483 352899 -1173 352915
rect -1483 352621 -1467 352899
rect -1189 352621 -1173 352899
rect -1483 334727 -1173 352621
rect -1483 334449 -1467 334727
rect -1189 334449 -1173 334727
rect -1483 316727 -1173 334449
rect -1483 316449 -1467 316727
rect -1189 316449 -1173 316727
rect -1483 298727 -1173 316449
rect -1483 298449 -1467 298727
rect -1189 298449 -1173 298727
rect -1483 280727 -1173 298449
rect -1483 280449 -1467 280727
rect -1189 280449 -1173 280727
rect -1483 262727 -1173 280449
rect -1483 262449 -1467 262727
rect -1189 262449 -1173 262727
rect -1483 244727 -1173 262449
rect -1483 244449 -1467 244727
rect -1189 244449 -1173 244727
rect -1483 226727 -1173 244449
rect -1483 226449 -1467 226727
rect -1189 226449 -1173 226727
rect -1483 208727 -1173 226449
rect -1483 208449 -1467 208727
rect -1189 208449 -1173 208727
rect -1483 190727 -1173 208449
rect -1483 190449 -1467 190727
rect -1189 190449 -1173 190727
rect -1483 172727 -1173 190449
rect -1483 172449 -1467 172727
rect -1189 172449 -1173 172727
rect -1483 154727 -1173 172449
rect -1483 154449 -1467 154727
rect -1189 154449 -1173 154727
rect -1483 136727 -1173 154449
rect -1483 136449 -1467 136727
rect -1189 136449 -1173 136727
rect -1483 118727 -1173 136449
rect -1483 118449 -1467 118727
rect -1189 118449 -1173 118727
rect -1483 100727 -1173 118449
rect -1483 100449 -1467 100727
rect -1189 100449 -1173 100727
rect -1483 82727 -1173 100449
rect -1483 82449 -1467 82727
rect -1189 82449 -1173 82727
rect -1483 64727 -1173 82449
rect -1483 64449 -1467 64727
rect -1189 64449 -1173 64727
rect -1483 46727 -1173 64449
rect -1483 46449 -1467 46727
rect -1189 46449 -1173 46727
rect -1483 28727 -1173 46449
rect -1483 28449 -1467 28727
rect -1189 28449 -1173 28727
rect -1483 10727 -1173 28449
rect -1483 10449 -1467 10727
rect -1189 10449 -1173 10727
rect -1483 -653 -1173 10449
rect -1003 352419 -693 352435
rect -1003 352141 -987 352419
rect -709 352141 -693 352419
rect -1003 343727 -693 352141
rect -1003 343449 -987 343727
rect -709 343449 -693 343727
rect -1003 325727 -693 343449
rect -1003 325449 -987 325727
rect -709 325449 -693 325727
rect -1003 307727 -693 325449
rect -1003 307449 -987 307727
rect -709 307449 -693 307727
rect -1003 289727 -693 307449
rect -1003 289449 -987 289727
rect -709 289449 -693 289727
rect -1003 271727 -693 289449
rect -1003 271449 -987 271727
rect -709 271449 -693 271727
rect -1003 253727 -693 271449
rect -1003 253449 -987 253727
rect -709 253449 -693 253727
rect -1003 235727 -693 253449
rect -1003 235449 -987 235727
rect -709 235449 -693 235727
rect -1003 217727 -693 235449
rect -1003 217449 -987 217727
rect -709 217449 -693 217727
rect -1003 199727 -693 217449
rect -1003 199449 -987 199727
rect -709 199449 -693 199727
rect -1003 181727 -693 199449
rect -1003 181449 -987 181727
rect -709 181449 -693 181727
rect -1003 163727 -693 181449
rect -1003 163449 -987 163727
rect -709 163449 -693 163727
rect -1003 145727 -693 163449
rect -1003 145449 -987 145727
rect -709 145449 -693 145727
rect -1003 127727 -693 145449
rect -1003 127449 -987 127727
rect -709 127449 -693 127727
rect -1003 109727 -693 127449
rect -1003 109449 -987 109727
rect -709 109449 -693 109727
rect -1003 91727 -693 109449
rect -1003 91449 -987 91727
rect -709 91449 -693 91727
rect -1003 73727 -693 91449
rect -1003 73449 -987 73727
rect -709 73449 -693 73727
rect -1003 55727 -693 73449
rect -1003 55449 -987 55727
rect -709 55449 -693 55727
rect -1003 37727 -693 55449
rect -1003 37449 -987 37727
rect -709 37449 -693 37727
rect -1003 19727 -693 37449
rect -1003 19449 -987 19727
rect -709 19449 -693 19727
rect -1003 1727 -693 19449
rect -1003 1449 -987 1727
rect -709 1449 -693 1727
rect -1003 -173 -693 1449
rect -1003 -451 -987 -173
rect -709 -451 -693 -173
rect -1003 -467 -693 -451
rect 897 352419 1207 352915
rect 897 352141 913 352419
rect 1191 352141 1207 352419
rect 897 343727 1207 352141
rect 897 343449 913 343727
rect 1191 343449 1207 343727
rect 897 325727 1207 343449
rect 897 325449 913 325727
rect 1191 325449 1207 325727
rect 897 307727 1207 325449
rect 897 307449 913 307727
rect 1191 307449 1207 307727
rect 897 289727 1207 307449
rect 897 289449 913 289727
rect 1191 289449 1207 289727
rect 897 271727 1207 289449
rect 897 271449 913 271727
rect 1191 271449 1207 271727
rect 897 253727 1207 271449
rect 897 253449 913 253727
rect 1191 253449 1207 253727
rect 897 235727 1207 253449
rect 897 235449 913 235727
rect 1191 235449 1207 235727
rect 897 217727 1207 235449
rect 897 217449 913 217727
rect 1191 217449 1207 217727
rect 897 199727 1207 217449
rect 897 199449 913 199727
rect 1191 199449 1207 199727
rect 897 181727 1207 199449
rect 897 181449 913 181727
rect 1191 181449 1207 181727
rect 897 163727 1207 181449
rect 897 163449 913 163727
rect 1191 163449 1207 163727
rect 897 145727 1207 163449
rect 897 145449 913 145727
rect 1191 145449 1207 145727
rect 897 127727 1207 145449
rect 897 127449 913 127727
rect 1191 127449 1207 127727
rect 897 109727 1207 127449
rect 897 109449 913 109727
rect 1191 109449 1207 109727
rect 897 91727 1207 109449
rect 897 91449 913 91727
rect 1191 91449 1207 91727
rect 897 73727 1207 91449
rect 897 73449 913 73727
rect 1191 73449 1207 73727
rect 897 55727 1207 73449
rect 897 55449 913 55727
rect 1191 55449 1207 55727
rect 897 37727 1207 55449
rect 897 37449 913 37727
rect 1191 37449 1207 37727
rect 897 19727 1207 37449
rect 897 19449 913 19727
rect 1191 19449 1207 19727
rect 897 1727 1207 19449
rect 897 1449 913 1727
rect 1191 1449 1207 1727
rect 897 -173 1207 1449
rect 897 -451 913 -173
rect 1191 -451 1207 -173
rect -1483 -931 -1467 -653
rect -1189 -931 -1173 -653
rect -1483 -947 -1173 -931
rect 897 -947 1207 -451
rect 2757 345587 3067 353101
rect 2757 345309 2773 345587
rect 3051 345309 3067 345587
rect 2757 327587 3067 345309
rect 2757 327309 2773 327587
rect 3051 327309 3067 327587
rect 2757 309587 3067 327309
rect 2757 309309 2773 309587
rect 3051 309309 3067 309587
rect 2757 291587 3067 309309
rect 2757 291309 2773 291587
rect 3051 291309 3067 291587
rect 2757 273587 3067 291309
rect 2757 273309 2773 273587
rect 3051 273309 3067 273587
rect 2757 255587 3067 273309
rect 2757 255309 2773 255587
rect 3051 255309 3067 255587
rect 2757 237587 3067 255309
rect 2757 237309 2773 237587
rect 3051 237309 3067 237587
rect 2757 219587 3067 237309
rect 2757 219309 2773 219587
rect 3051 219309 3067 219587
rect 2757 201587 3067 219309
rect 2757 201309 2773 201587
rect 3051 201309 3067 201587
rect 2757 183587 3067 201309
rect 2757 183309 2773 183587
rect 3051 183309 3067 183587
rect 2757 165587 3067 183309
rect 2757 165309 2773 165587
rect 3051 165309 3067 165587
rect 2757 147587 3067 165309
rect 2757 147309 2773 147587
rect 3051 147309 3067 147587
rect 2757 129587 3067 147309
rect 2757 129309 2773 129587
rect 3051 129309 3067 129587
rect 2757 111587 3067 129309
rect 2757 111309 2773 111587
rect 3051 111309 3067 111587
rect 2757 93587 3067 111309
rect 2757 93309 2773 93587
rect 3051 93309 3067 93587
rect 2757 75587 3067 93309
rect 2757 75309 2773 75587
rect 3051 75309 3067 75587
rect 2757 57587 3067 75309
rect 2757 57309 2773 57587
rect 3051 57309 3067 57587
rect 2757 39587 3067 57309
rect 2757 39309 2773 39587
rect 3051 39309 3067 39587
rect 2757 21587 3067 39309
rect 2757 21309 2773 21587
rect 3051 21309 3067 21587
rect 2757 3587 3067 21309
rect 2757 3309 2773 3587
rect 3051 3309 3067 3587
rect -1963 -1411 -1947 -1133
rect -1669 -1411 -1653 -1133
rect -1963 -1427 -1653 -1411
rect 2757 -1133 3067 3309
rect 2757 -1411 2773 -1133
rect 3051 -1411 3067 -1133
rect -2443 -1891 -2427 -1613
rect -2149 -1891 -2133 -1613
rect -2443 -1907 -2133 -1891
rect 2757 -1907 3067 -1411
rect 4617 347447 4927 354061
rect 4617 347169 4633 347447
rect 4911 347169 4927 347447
rect 4617 329447 4927 347169
rect 4617 329169 4633 329447
rect 4911 329169 4927 329447
rect 4617 311447 4927 329169
rect 4617 311169 4633 311447
rect 4911 311169 4927 311447
rect 4617 293447 4927 311169
rect 4617 293169 4633 293447
rect 4911 293169 4927 293447
rect 4617 275447 4927 293169
rect 4617 275169 4633 275447
rect 4911 275169 4927 275447
rect 4617 257447 4927 275169
rect 4617 257169 4633 257447
rect 4911 257169 4927 257447
rect 4617 239447 4927 257169
rect 4617 239169 4633 239447
rect 4911 239169 4927 239447
rect 4617 221447 4927 239169
rect 4617 221169 4633 221447
rect 4911 221169 4927 221447
rect 4617 203447 4927 221169
rect 4617 203169 4633 203447
rect 4911 203169 4927 203447
rect 4617 185447 4927 203169
rect 4617 185169 4633 185447
rect 4911 185169 4927 185447
rect 4617 167447 4927 185169
rect 4617 167169 4633 167447
rect 4911 167169 4927 167447
rect 4617 149447 4927 167169
rect 4617 149169 4633 149447
rect 4911 149169 4927 149447
rect 4617 131447 4927 149169
rect 4617 131169 4633 131447
rect 4911 131169 4927 131447
rect 4617 113447 4927 131169
rect 4617 113169 4633 113447
rect 4911 113169 4927 113447
rect 4617 95447 4927 113169
rect 4617 95169 4633 95447
rect 4911 95169 4927 95447
rect 4617 77447 4927 95169
rect 4617 77169 4633 77447
rect 4911 77169 4927 77447
rect 4617 59447 4927 77169
rect 4617 59169 4633 59447
rect 4911 59169 4927 59447
rect 4617 41447 4927 59169
rect 4617 41169 4633 41447
rect 4911 41169 4927 41447
rect 4617 23447 4927 41169
rect 4617 23169 4633 23447
rect 4911 23169 4927 23447
rect 4617 5447 4927 23169
rect 4617 5169 4633 5447
rect 4911 5169 4927 5447
rect -2923 -2371 -2907 -2093
rect -2629 -2371 -2613 -2093
rect -2923 -2387 -2613 -2371
rect 4617 -2093 4927 5169
rect 4617 -2371 4633 -2093
rect 4911 -2371 4927 -2093
rect -3403 -2851 -3387 -2573
rect -3109 -2851 -3093 -2573
rect -3403 -2867 -3093 -2851
rect 4617 -2867 4927 -2371
rect 6477 349307 6787 355021
rect 15477 355779 15787 355795
rect 15477 355501 15493 355779
rect 15771 355501 15787 355779
rect 13617 354819 13927 354835
rect 13617 354541 13633 354819
rect 13911 354541 13927 354819
rect 11757 353859 12067 353875
rect 11757 353581 11773 353859
rect 12051 353581 12067 353859
rect 6477 349029 6493 349307
rect 6771 349029 6787 349307
rect 6477 331307 6787 349029
rect 6477 331029 6493 331307
rect 6771 331029 6787 331307
rect 6477 313307 6787 331029
rect 6477 313029 6493 313307
rect 6771 313029 6787 313307
rect 6477 295307 6787 313029
rect 6477 295029 6493 295307
rect 6771 295029 6787 295307
rect 6477 277307 6787 295029
rect 6477 277029 6493 277307
rect 6771 277029 6787 277307
rect 6477 259307 6787 277029
rect 6477 259029 6493 259307
rect 6771 259029 6787 259307
rect 6477 241307 6787 259029
rect 6477 241029 6493 241307
rect 6771 241029 6787 241307
rect 6477 223307 6787 241029
rect 6477 223029 6493 223307
rect 6771 223029 6787 223307
rect 6477 205307 6787 223029
rect 6477 205029 6493 205307
rect 6771 205029 6787 205307
rect 6477 187307 6787 205029
rect 6477 187029 6493 187307
rect 6771 187029 6787 187307
rect 6477 169307 6787 187029
rect 6477 169029 6493 169307
rect 6771 169029 6787 169307
rect 6477 151307 6787 169029
rect 6477 151029 6493 151307
rect 6771 151029 6787 151307
rect 6477 133307 6787 151029
rect 6477 133029 6493 133307
rect 6771 133029 6787 133307
rect 6477 115307 6787 133029
rect 6477 115029 6493 115307
rect 6771 115029 6787 115307
rect 6477 97307 6787 115029
rect 6477 97029 6493 97307
rect 6771 97029 6787 97307
rect 6477 79307 6787 97029
rect 6477 79029 6493 79307
rect 6771 79029 6787 79307
rect 6477 61307 6787 79029
rect 6477 61029 6493 61307
rect 6771 61029 6787 61307
rect 6477 43307 6787 61029
rect 6477 43029 6493 43307
rect 6771 43029 6787 43307
rect 6477 25307 6787 43029
rect 6477 25029 6493 25307
rect 6771 25029 6787 25307
rect 6477 7307 6787 25029
rect 6477 7029 6493 7307
rect 6771 7029 6787 7307
rect -3883 -3331 -3867 -3053
rect -3589 -3331 -3573 -3053
rect -3883 -3347 -3573 -3331
rect 6477 -3053 6787 7029
rect 9897 352899 10207 352915
rect 9897 352621 9913 352899
rect 10191 352621 10207 352899
rect 9897 334727 10207 352621
rect 9897 334449 9913 334727
rect 10191 334449 10207 334727
rect 9897 316727 10207 334449
rect 9897 316449 9913 316727
rect 10191 316449 10207 316727
rect 9897 298727 10207 316449
rect 9897 298449 9913 298727
rect 10191 298449 10207 298727
rect 9897 280727 10207 298449
rect 9897 280449 9913 280727
rect 10191 280449 10207 280727
rect 9897 262727 10207 280449
rect 9897 262449 9913 262727
rect 10191 262449 10207 262727
rect 9897 244727 10207 262449
rect 9897 244449 9913 244727
rect 10191 244449 10207 244727
rect 9897 226727 10207 244449
rect 9897 226449 9913 226727
rect 10191 226449 10207 226727
rect 9897 208727 10207 226449
rect 9897 208449 9913 208727
rect 10191 208449 10207 208727
rect 9897 190727 10207 208449
rect 9897 190449 9913 190727
rect 10191 190449 10207 190727
rect 9897 172727 10207 190449
rect 9897 172449 9913 172727
rect 10191 172449 10207 172727
rect 9897 154727 10207 172449
rect 9897 154449 9913 154727
rect 10191 154449 10207 154727
rect 9897 136727 10207 154449
rect 9897 136449 9913 136727
rect 10191 136449 10207 136727
rect 9897 118727 10207 136449
rect 9897 118449 9913 118727
rect 10191 118449 10207 118727
rect 9897 100727 10207 118449
rect 9897 100449 9913 100727
rect 10191 100449 10207 100727
rect 9897 82727 10207 100449
rect 9897 82449 9913 82727
rect 10191 82449 10207 82727
rect 9897 64727 10207 82449
rect 9897 64449 9913 64727
rect 10191 64449 10207 64727
rect 9897 46727 10207 64449
rect 9897 46449 9913 46727
rect 10191 46449 10207 46727
rect 9897 28727 10207 46449
rect 9897 28449 9913 28727
rect 10191 28449 10207 28727
rect 9897 10727 10207 28449
rect 9897 10449 9913 10727
rect 10191 10449 10207 10727
rect 9897 -653 10207 10449
rect 9897 -931 9913 -653
rect 10191 -931 10207 -653
rect 9897 -947 10207 -931
rect 11757 336587 12067 353581
rect 11757 336309 11773 336587
rect 12051 336309 12067 336587
rect 11757 318587 12067 336309
rect 11757 318309 11773 318587
rect 12051 318309 12067 318587
rect 11757 300587 12067 318309
rect 11757 300309 11773 300587
rect 12051 300309 12067 300587
rect 11757 282587 12067 300309
rect 11757 282309 11773 282587
rect 12051 282309 12067 282587
rect 11757 264587 12067 282309
rect 11757 264309 11773 264587
rect 12051 264309 12067 264587
rect 11757 246587 12067 264309
rect 11757 246309 11773 246587
rect 12051 246309 12067 246587
rect 11757 228587 12067 246309
rect 11757 228309 11773 228587
rect 12051 228309 12067 228587
rect 11757 210587 12067 228309
rect 11757 210309 11773 210587
rect 12051 210309 12067 210587
rect 11757 192587 12067 210309
rect 11757 192309 11773 192587
rect 12051 192309 12067 192587
rect 11757 174587 12067 192309
rect 11757 174309 11773 174587
rect 12051 174309 12067 174587
rect 11757 156587 12067 174309
rect 11757 156309 11773 156587
rect 12051 156309 12067 156587
rect 11757 138587 12067 156309
rect 11757 138309 11773 138587
rect 12051 138309 12067 138587
rect 11757 120587 12067 138309
rect 11757 120309 11773 120587
rect 12051 120309 12067 120587
rect 11757 102587 12067 120309
rect 11757 102309 11773 102587
rect 12051 102309 12067 102587
rect 11757 84587 12067 102309
rect 11757 84309 11773 84587
rect 12051 84309 12067 84587
rect 11757 66587 12067 84309
rect 11757 66309 11773 66587
rect 12051 66309 12067 66587
rect 11757 48587 12067 66309
rect 11757 48309 11773 48587
rect 12051 48309 12067 48587
rect 11757 30587 12067 48309
rect 11757 30309 11773 30587
rect 12051 30309 12067 30587
rect 11757 12587 12067 30309
rect 11757 12309 11773 12587
rect 12051 12309 12067 12587
rect 11757 -1613 12067 12309
rect 11757 -1891 11773 -1613
rect 12051 -1891 12067 -1613
rect 11757 -1907 12067 -1891
rect 13617 338447 13927 354541
rect 13617 338169 13633 338447
rect 13911 338169 13927 338447
rect 13617 320447 13927 338169
rect 13617 320169 13633 320447
rect 13911 320169 13927 320447
rect 13617 302447 13927 320169
rect 13617 302169 13633 302447
rect 13911 302169 13927 302447
rect 13617 284447 13927 302169
rect 13617 284169 13633 284447
rect 13911 284169 13927 284447
rect 13617 266447 13927 284169
rect 13617 266169 13633 266447
rect 13911 266169 13927 266447
rect 13617 248447 13927 266169
rect 13617 248169 13633 248447
rect 13911 248169 13927 248447
rect 13617 230447 13927 248169
rect 13617 230169 13633 230447
rect 13911 230169 13927 230447
rect 13617 212447 13927 230169
rect 13617 212169 13633 212447
rect 13911 212169 13927 212447
rect 13617 194447 13927 212169
rect 13617 194169 13633 194447
rect 13911 194169 13927 194447
rect 13617 176447 13927 194169
rect 13617 176169 13633 176447
rect 13911 176169 13927 176447
rect 13617 158447 13927 176169
rect 13617 158169 13633 158447
rect 13911 158169 13927 158447
rect 13617 140447 13927 158169
rect 13617 140169 13633 140447
rect 13911 140169 13927 140447
rect 13617 122447 13927 140169
rect 13617 122169 13633 122447
rect 13911 122169 13927 122447
rect 13617 104447 13927 122169
rect 13617 104169 13633 104447
rect 13911 104169 13927 104447
rect 13617 86447 13927 104169
rect 13617 86169 13633 86447
rect 13911 86169 13927 86447
rect 13617 68447 13927 86169
rect 13617 68169 13633 68447
rect 13911 68169 13927 68447
rect 13617 50447 13927 68169
rect 13617 50169 13633 50447
rect 13911 50169 13927 50447
rect 13617 32447 13927 50169
rect 13617 32169 13633 32447
rect 13911 32169 13927 32447
rect 13617 14447 13927 32169
rect 13617 14169 13633 14447
rect 13911 14169 13927 14447
rect 13617 -2573 13927 14169
rect 13617 -2851 13633 -2573
rect 13911 -2851 13927 -2573
rect 13617 -2867 13927 -2851
rect 15477 340307 15787 355501
rect 24477 355299 24787 355795
rect 24477 355021 24493 355299
rect 24771 355021 24787 355299
rect 22617 354339 22927 354835
rect 22617 354061 22633 354339
rect 22911 354061 22927 354339
rect 20757 353379 21067 353875
rect 20757 353101 20773 353379
rect 21051 353101 21067 353379
rect 15477 340029 15493 340307
rect 15771 340029 15787 340307
rect 15477 322307 15787 340029
rect 15477 322029 15493 322307
rect 15771 322029 15787 322307
rect 15477 304307 15787 322029
rect 15477 304029 15493 304307
rect 15771 304029 15787 304307
rect 15477 286307 15787 304029
rect 15477 286029 15493 286307
rect 15771 286029 15787 286307
rect 15477 268307 15787 286029
rect 15477 268029 15493 268307
rect 15771 268029 15787 268307
rect 15477 250307 15787 268029
rect 15477 250029 15493 250307
rect 15771 250029 15787 250307
rect 15477 232307 15787 250029
rect 15477 232029 15493 232307
rect 15771 232029 15787 232307
rect 15477 214307 15787 232029
rect 15477 214029 15493 214307
rect 15771 214029 15787 214307
rect 15477 196307 15787 214029
rect 15477 196029 15493 196307
rect 15771 196029 15787 196307
rect 15477 178307 15787 196029
rect 15477 178029 15493 178307
rect 15771 178029 15787 178307
rect 15477 160307 15787 178029
rect 15477 160029 15493 160307
rect 15771 160029 15787 160307
rect 15477 142307 15787 160029
rect 15477 142029 15493 142307
rect 15771 142029 15787 142307
rect 15477 124307 15787 142029
rect 15477 124029 15493 124307
rect 15771 124029 15787 124307
rect 15477 106307 15787 124029
rect 15477 106029 15493 106307
rect 15771 106029 15787 106307
rect 15477 88307 15787 106029
rect 15477 88029 15493 88307
rect 15771 88029 15787 88307
rect 15477 70307 15787 88029
rect 15477 70029 15493 70307
rect 15771 70029 15787 70307
rect 15477 52307 15787 70029
rect 15477 52029 15493 52307
rect 15771 52029 15787 52307
rect 15477 34307 15787 52029
rect 15477 34029 15493 34307
rect 15771 34029 15787 34307
rect 15477 16307 15787 34029
rect 15477 16029 15493 16307
rect 15771 16029 15787 16307
rect 6477 -3331 6493 -3053
rect 6771 -3331 6787 -3053
rect -4363 -3811 -4347 -3533
rect -4069 -3811 -4053 -3533
rect -4363 -3827 -4053 -3811
rect 6477 -3827 6787 -3331
rect 15477 -3533 15787 16029
rect 18897 352419 19207 352915
rect 18897 352141 18913 352419
rect 19191 352141 19207 352419
rect 18897 343727 19207 352141
rect 18897 343449 18913 343727
rect 19191 343449 19207 343727
rect 18897 325727 19207 343449
rect 18897 325449 18913 325727
rect 19191 325449 19207 325727
rect 18897 307727 19207 325449
rect 18897 307449 18913 307727
rect 19191 307449 19207 307727
rect 18897 289727 19207 307449
rect 18897 289449 18913 289727
rect 19191 289449 19207 289727
rect 18897 271727 19207 289449
rect 18897 271449 18913 271727
rect 19191 271449 19207 271727
rect 18897 253727 19207 271449
rect 18897 253449 18913 253727
rect 19191 253449 19207 253727
rect 18897 235727 19207 253449
rect 18897 235449 18913 235727
rect 19191 235449 19207 235727
rect 18897 217727 19207 235449
rect 18897 217449 18913 217727
rect 19191 217449 19207 217727
rect 18897 199727 19207 217449
rect 18897 199449 18913 199727
rect 19191 199449 19207 199727
rect 18897 181727 19207 199449
rect 18897 181449 18913 181727
rect 19191 181449 19207 181727
rect 18897 163727 19207 181449
rect 18897 163449 18913 163727
rect 19191 163449 19207 163727
rect 18897 145727 19207 163449
rect 18897 145449 18913 145727
rect 19191 145449 19207 145727
rect 18897 127727 19207 145449
rect 18897 127449 18913 127727
rect 19191 127449 19207 127727
rect 18897 109727 19207 127449
rect 18897 109449 18913 109727
rect 19191 109449 19207 109727
rect 18897 91727 19207 109449
rect 18897 91449 18913 91727
rect 19191 91449 19207 91727
rect 18897 73727 19207 91449
rect 18897 73449 18913 73727
rect 19191 73449 19207 73727
rect 18897 55727 19207 73449
rect 18897 55449 18913 55727
rect 19191 55449 19207 55727
rect 18897 37727 19207 55449
rect 18897 37449 18913 37727
rect 19191 37449 19207 37727
rect 18897 19727 19207 37449
rect 18897 19449 18913 19727
rect 19191 19449 19207 19727
rect 18897 1727 19207 19449
rect 18897 1449 18913 1727
rect 19191 1449 19207 1727
rect 18897 -173 19207 1449
rect 18897 -451 18913 -173
rect 19191 -451 19207 -173
rect 18897 -947 19207 -451
rect 20757 345587 21067 353101
rect 20757 345309 20773 345587
rect 21051 345309 21067 345587
rect 20757 327587 21067 345309
rect 20757 327309 20773 327587
rect 21051 327309 21067 327587
rect 20757 309587 21067 327309
rect 20757 309309 20773 309587
rect 21051 309309 21067 309587
rect 20757 291587 21067 309309
rect 20757 291309 20773 291587
rect 21051 291309 21067 291587
rect 20757 273587 21067 291309
rect 20757 273309 20773 273587
rect 21051 273309 21067 273587
rect 20757 255587 21067 273309
rect 20757 255309 20773 255587
rect 21051 255309 21067 255587
rect 20757 237587 21067 255309
rect 20757 237309 20773 237587
rect 21051 237309 21067 237587
rect 20757 219587 21067 237309
rect 20757 219309 20773 219587
rect 21051 219309 21067 219587
rect 20757 201587 21067 219309
rect 20757 201309 20773 201587
rect 21051 201309 21067 201587
rect 20757 183587 21067 201309
rect 20757 183309 20773 183587
rect 21051 183309 21067 183587
rect 20757 165587 21067 183309
rect 20757 165309 20773 165587
rect 21051 165309 21067 165587
rect 20757 147587 21067 165309
rect 20757 147309 20773 147587
rect 21051 147309 21067 147587
rect 20757 129587 21067 147309
rect 20757 129309 20773 129587
rect 21051 129309 21067 129587
rect 20757 111587 21067 129309
rect 20757 111309 20773 111587
rect 21051 111309 21067 111587
rect 20757 93587 21067 111309
rect 20757 93309 20773 93587
rect 21051 93309 21067 93587
rect 20757 75587 21067 93309
rect 20757 75309 20773 75587
rect 21051 75309 21067 75587
rect 20757 57587 21067 75309
rect 20757 57309 20773 57587
rect 21051 57309 21067 57587
rect 20757 39587 21067 57309
rect 20757 39309 20773 39587
rect 21051 39309 21067 39587
rect 20757 21587 21067 39309
rect 20757 21309 20773 21587
rect 21051 21309 21067 21587
rect 20757 3587 21067 21309
rect 20757 3309 20773 3587
rect 21051 3309 21067 3587
rect 20757 -1133 21067 3309
rect 20757 -1411 20773 -1133
rect 21051 -1411 21067 -1133
rect 20757 -1907 21067 -1411
rect 22617 347447 22927 354061
rect 22617 347169 22633 347447
rect 22911 347169 22927 347447
rect 22617 329447 22927 347169
rect 22617 329169 22633 329447
rect 22911 329169 22927 329447
rect 22617 311447 22927 329169
rect 22617 311169 22633 311447
rect 22911 311169 22927 311447
rect 22617 293447 22927 311169
rect 22617 293169 22633 293447
rect 22911 293169 22927 293447
rect 22617 275447 22927 293169
rect 22617 275169 22633 275447
rect 22911 275169 22927 275447
rect 22617 257447 22927 275169
rect 22617 257169 22633 257447
rect 22911 257169 22927 257447
rect 22617 239447 22927 257169
rect 22617 239169 22633 239447
rect 22911 239169 22927 239447
rect 22617 221447 22927 239169
rect 22617 221169 22633 221447
rect 22911 221169 22927 221447
rect 22617 203447 22927 221169
rect 22617 203169 22633 203447
rect 22911 203169 22927 203447
rect 22617 185447 22927 203169
rect 22617 185169 22633 185447
rect 22911 185169 22927 185447
rect 22617 167447 22927 185169
rect 22617 167169 22633 167447
rect 22911 167169 22927 167447
rect 22617 149447 22927 167169
rect 22617 149169 22633 149447
rect 22911 149169 22927 149447
rect 22617 131447 22927 149169
rect 22617 131169 22633 131447
rect 22911 131169 22927 131447
rect 22617 113447 22927 131169
rect 22617 113169 22633 113447
rect 22911 113169 22927 113447
rect 22617 95447 22927 113169
rect 22617 95169 22633 95447
rect 22911 95169 22927 95447
rect 22617 77447 22927 95169
rect 22617 77169 22633 77447
rect 22911 77169 22927 77447
rect 22617 59447 22927 77169
rect 22617 59169 22633 59447
rect 22911 59169 22927 59447
rect 22617 41447 22927 59169
rect 22617 41169 22633 41447
rect 22911 41169 22927 41447
rect 22617 23447 22927 41169
rect 22617 23169 22633 23447
rect 22911 23169 22927 23447
rect 22617 5447 22927 23169
rect 22617 5169 22633 5447
rect 22911 5169 22927 5447
rect 22617 -2093 22927 5169
rect 22617 -2371 22633 -2093
rect 22911 -2371 22927 -2093
rect 22617 -2867 22927 -2371
rect 24477 349307 24787 355021
rect 33477 355779 33787 355795
rect 33477 355501 33493 355779
rect 33771 355501 33787 355779
rect 31617 354819 31927 354835
rect 31617 354541 31633 354819
rect 31911 354541 31927 354819
rect 29757 353859 30067 353875
rect 29757 353581 29773 353859
rect 30051 353581 30067 353859
rect 24477 349029 24493 349307
rect 24771 349029 24787 349307
rect 24477 331307 24787 349029
rect 24477 331029 24493 331307
rect 24771 331029 24787 331307
rect 24477 313307 24787 331029
rect 24477 313029 24493 313307
rect 24771 313029 24787 313307
rect 24477 295307 24787 313029
rect 24477 295029 24493 295307
rect 24771 295029 24787 295307
rect 24477 277307 24787 295029
rect 24477 277029 24493 277307
rect 24771 277029 24787 277307
rect 24477 259307 24787 277029
rect 24477 259029 24493 259307
rect 24771 259029 24787 259307
rect 24477 241307 24787 259029
rect 24477 241029 24493 241307
rect 24771 241029 24787 241307
rect 24477 223307 24787 241029
rect 24477 223029 24493 223307
rect 24771 223029 24787 223307
rect 24477 205307 24787 223029
rect 24477 205029 24493 205307
rect 24771 205029 24787 205307
rect 24477 187307 24787 205029
rect 24477 187029 24493 187307
rect 24771 187029 24787 187307
rect 24477 169307 24787 187029
rect 24477 169029 24493 169307
rect 24771 169029 24787 169307
rect 24477 151307 24787 169029
rect 24477 151029 24493 151307
rect 24771 151029 24787 151307
rect 24477 133307 24787 151029
rect 24477 133029 24493 133307
rect 24771 133029 24787 133307
rect 24477 115307 24787 133029
rect 24477 115029 24493 115307
rect 24771 115029 24787 115307
rect 24477 97307 24787 115029
rect 24477 97029 24493 97307
rect 24771 97029 24787 97307
rect 24477 79307 24787 97029
rect 24477 79029 24493 79307
rect 24771 79029 24787 79307
rect 24477 61307 24787 79029
rect 24477 61029 24493 61307
rect 24771 61029 24787 61307
rect 24477 43307 24787 61029
rect 24477 43029 24493 43307
rect 24771 43029 24787 43307
rect 24477 25307 24787 43029
rect 24477 25029 24493 25307
rect 24771 25029 24787 25307
rect 24477 7307 24787 25029
rect 24477 7029 24493 7307
rect 24771 7029 24787 7307
rect 15477 -3811 15493 -3533
rect 15771 -3811 15787 -3533
rect 15477 -3827 15787 -3811
rect 24477 -3053 24787 7029
rect 27897 352899 28207 352915
rect 27897 352621 27913 352899
rect 28191 352621 28207 352899
rect 27897 334727 28207 352621
rect 27897 334449 27913 334727
rect 28191 334449 28207 334727
rect 27897 316727 28207 334449
rect 27897 316449 27913 316727
rect 28191 316449 28207 316727
rect 27897 298727 28207 316449
rect 27897 298449 27913 298727
rect 28191 298449 28207 298727
rect 27897 280727 28207 298449
rect 27897 280449 27913 280727
rect 28191 280449 28207 280727
rect 27897 262727 28207 280449
rect 27897 262449 27913 262727
rect 28191 262449 28207 262727
rect 27897 244727 28207 262449
rect 27897 244449 27913 244727
rect 28191 244449 28207 244727
rect 27897 226727 28207 244449
rect 27897 226449 27913 226727
rect 28191 226449 28207 226727
rect 27897 208727 28207 226449
rect 27897 208449 27913 208727
rect 28191 208449 28207 208727
rect 27897 190727 28207 208449
rect 27897 190449 27913 190727
rect 28191 190449 28207 190727
rect 27897 172727 28207 190449
rect 27897 172449 27913 172727
rect 28191 172449 28207 172727
rect 27897 154727 28207 172449
rect 27897 154449 27913 154727
rect 28191 154449 28207 154727
rect 27897 136727 28207 154449
rect 27897 136449 27913 136727
rect 28191 136449 28207 136727
rect 27897 118727 28207 136449
rect 27897 118449 27913 118727
rect 28191 118449 28207 118727
rect 27897 100727 28207 118449
rect 27897 100449 27913 100727
rect 28191 100449 28207 100727
rect 27897 82727 28207 100449
rect 27897 82449 27913 82727
rect 28191 82449 28207 82727
rect 27897 64727 28207 82449
rect 27897 64449 27913 64727
rect 28191 64449 28207 64727
rect 27897 46727 28207 64449
rect 27897 46449 27913 46727
rect 28191 46449 28207 46727
rect 27897 28727 28207 46449
rect 27897 28449 27913 28727
rect 28191 28449 28207 28727
rect 27897 10727 28207 28449
rect 27897 10449 27913 10727
rect 28191 10449 28207 10727
rect 27897 -653 28207 10449
rect 27897 -931 27913 -653
rect 28191 -931 28207 -653
rect 27897 -947 28207 -931
rect 29757 336587 30067 353581
rect 29757 336309 29773 336587
rect 30051 336309 30067 336587
rect 29757 318587 30067 336309
rect 29757 318309 29773 318587
rect 30051 318309 30067 318587
rect 29757 300587 30067 318309
rect 29757 300309 29773 300587
rect 30051 300309 30067 300587
rect 29757 282587 30067 300309
rect 29757 282309 29773 282587
rect 30051 282309 30067 282587
rect 29757 264587 30067 282309
rect 29757 264309 29773 264587
rect 30051 264309 30067 264587
rect 29757 246587 30067 264309
rect 29757 246309 29773 246587
rect 30051 246309 30067 246587
rect 29757 228587 30067 246309
rect 29757 228309 29773 228587
rect 30051 228309 30067 228587
rect 29757 210587 30067 228309
rect 29757 210309 29773 210587
rect 30051 210309 30067 210587
rect 29757 192587 30067 210309
rect 29757 192309 29773 192587
rect 30051 192309 30067 192587
rect 29757 174587 30067 192309
rect 29757 174309 29773 174587
rect 30051 174309 30067 174587
rect 29757 156587 30067 174309
rect 29757 156309 29773 156587
rect 30051 156309 30067 156587
rect 29757 138587 30067 156309
rect 29757 138309 29773 138587
rect 30051 138309 30067 138587
rect 29757 120587 30067 138309
rect 29757 120309 29773 120587
rect 30051 120309 30067 120587
rect 29757 102587 30067 120309
rect 29757 102309 29773 102587
rect 30051 102309 30067 102587
rect 29757 84587 30067 102309
rect 29757 84309 29773 84587
rect 30051 84309 30067 84587
rect 29757 66587 30067 84309
rect 29757 66309 29773 66587
rect 30051 66309 30067 66587
rect 29757 48587 30067 66309
rect 29757 48309 29773 48587
rect 30051 48309 30067 48587
rect 29757 30587 30067 48309
rect 29757 30309 29773 30587
rect 30051 30309 30067 30587
rect 29757 12587 30067 30309
rect 29757 12309 29773 12587
rect 30051 12309 30067 12587
rect 29757 -1613 30067 12309
rect 29757 -1891 29773 -1613
rect 30051 -1891 30067 -1613
rect 29757 -1907 30067 -1891
rect 31617 338447 31927 354541
rect 31617 338169 31633 338447
rect 31911 338169 31927 338447
rect 31617 320447 31927 338169
rect 31617 320169 31633 320447
rect 31911 320169 31927 320447
rect 31617 302447 31927 320169
rect 31617 302169 31633 302447
rect 31911 302169 31927 302447
rect 31617 284447 31927 302169
rect 31617 284169 31633 284447
rect 31911 284169 31927 284447
rect 31617 266447 31927 284169
rect 31617 266169 31633 266447
rect 31911 266169 31927 266447
rect 31617 248447 31927 266169
rect 31617 248169 31633 248447
rect 31911 248169 31927 248447
rect 31617 230447 31927 248169
rect 31617 230169 31633 230447
rect 31911 230169 31927 230447
rect 31617 212447 31927 230169
rect 31617 212169 31633 212447
rect 31911 212169 31927 212447
rect 31617 194447 31927 212169
rect 31617 194169 31633 194447
rect 31911 194169 31927 194447
rect 31617 176447 31927 194169
rect 31617 176169 31633 176447
rect 31911 176169 31927 176447
rect 31617 158447 31927 176169
rect 31617 158169 31633 158447
rect 31911 158169 31927 158447
rect 31617 140447 31927 158169
rect 31617 140169 31633 140447
rect 31911 140169 31927 140447
rect 31617 122447 31927 140169
rect 31617 122169 31633 122447
rect 31911 122169 31927 122447
rect 31617 104447 31927 122169
rect 31617 104169 31633 104447
rect 31911 104169 31927 104447
rect 31617 86447 31927 104169
rect 31617 86169 31633 86447
rect 31911 86169 31927 86447
rect 31617 68447 31927 86169
rect 31617 68169 31633 68447
rect 31911 68169 31927 68447
rect 31617 50447 31927 68169
rect 31617 50169 31633 50447
rect 31911 50169 31927 50447
rect 31617 32447 31927 50169
rect 31617 32169 31633 32447
rect 31911 32169 31927 32447
rect 31617 14447 31927 32169
rect 31617 14169 31633 14447
rect 31911 14169 31927 14447
rect 31617 -2573 31927 14169
rect 31617 -2851 31633 -2573
rect 31911 -2851 31927 -2573
rect 31617 -2867 31927 -2851
rect 33477 340307 33787 355501
rect 42477 355299 42787 355795
rect 42477 355021 42493 355299
rect 42771 355021 42787 355299
rect 40617 354339 40927 354835
rect 40617 354061 40633 354339
rect 40911 354061 40927 354339
rect 38757 353379 39067 353875
rect 38757 353101 38773 353379
rect 39051 353101 39067 353379
rect 33477 340029 33493 340307
rect 33771 340029 33787 340307
rect 33477 322307 33787 340029
rect 33477 322029 33493 322307
rect 33771 322029 33787 322307
rect 33477 304307 33787 322029
rect 33477 304029 33493 304307
rect 33771 304029 33787 304307
rect 33477 286307 33787 304029
rect 33477 286029 33493 286307
rect 33771 286029 33787 286307
rect 33477 268307 33787 286029
rect 33477 268029 33493 268307
rect 33771 268029 33787 268307
rect 33477 250307 33787 268029
rect 33477 250029 33493 250307
rect 33771 250029 33787 250307
rect 33477 232307 33787 250029
rect 33477 232029 33493 232307
rect 33771 232029 33787 232307
rect 33477 214307 33787 232029
rect 33477 214029 33493 214307
rect 33771 214029 33787 214307
rect 33477 196307 33787 214029
rect 33477 196029 33493 196307
rect 33771 196029 33787 196307
rect 33477 178307 33787 196029
rect 33477 178029 33493 178307
rect 33771 178029 33787 178307
rect 33477 160307 33787 178029
rect 33477 160029 33493 160307
rect 33771 160029 33787 160307
rect 33477 142307 33787 160029
rect 33477 142029 33493 142307
rect 33771 142029 33787 142307
rect 33477 124307 33787 142029
rect 33477 124029 33493 124307
rect 33771 124029 33787 124307
rect 33477 106307 33787 124029
rect 33477 106029 33493 106307
rect 33771 106029 33787 106307
rect 33477 88307 33787 106029
rect 33477 88029 33493 88307
rect 33771 88029 33787 88307
rect 33477 70307 33787 88029
rect 33477 70029 33493 70307
rect 33771 70029 33787 70307
rect 33477 52307 33787 70029
rect 33477 52029 33493 52307
rect 33771 52029 33787 52307
rect 33477 34307 33787 52029
rect 33477 34029 33493 34307
rect 33771 34029 33787 34307
rect 33477 16307 33787 34029
rect 33477 16029 33493 16307
rect 33771 16029 33787 16307
rect 24477 -3331 24493 -3053
rect 24771 -3331 24787 -3053
rect 24477 -3827 24787 -3331
rect 33477 -3533 33787 16029
rect 36897 352419 37207 352915
rect 36897 352141 36913 352419
rect 37191 352141 37207 352419
rect 36897 343727 37207 352141
rect 36897 343449 36913 343727
rect 37191 343449 37207 343727
rect 36897 325727 37207 343449
rect 36897 325449 36913 325727
rect 37191 325449 37207 325727
rect 36897 307727 37207 325449
rect 36897 307449 36913 307727
rect 37191 307449 37207 307727
rect 36897 289727 37207 307449
rect 36897 289449 36913 289727
rect 37191 289449 37207 289727
rect 36897 271727 37207 289449
rect 36897 271449 36913 271727
rect 37191 271449 37207 271727
rect 36897 253727 37207 271449
rect 36897 253449 36913 253727
rect 37191 253449 37207 253727
rect 36897 235727 37207 253449
rect 36897 235449 36913 235727
rect 37191 235449 37207 235727
rect 36897 217727 37207 235449
rect 36897 217449 36913 217727
rect 37191 217449 37207 217727
rect 36897 199727 37207 217449
rect 36897 199449 36913 199727
rect 37191 199449 37207 199727
rect 36897 181727 37207 199449
rect 36897 181449 36913 181727
rect 37191 181449 37207 181727
rect 36897 163727 37207 181449
rect 36897 163449 36913 163727
rect 37191 163449 37207 163727
rect 36897 145727 37207 163449
rect 36897 145449 36913 145727
rect 37191 145449 37207 145727
rect 36897 127727 37207 145449
rect 36897 127449 36913 127727
rect 37191 127449 37207 127727
rect 36897 109727 37207 127449
rect 36897 109449 36913 109727
rect 37191 109449 37207 109727
rect 36897 91727 37207 109449
rect 36897 91449 36913 91727
rect 37191 91449 37207 91727
rect 36897 73727 37207 91449
rect 36897 73449 36913 73727
rect 37191 73449 37207 73727
rect 36897 55727 37207 73449
rect 36897 55449 36913 55727
rect 37191 55449 37207 55727
rect 36897 37727 37207 55449
rect 36897 37449 36913 37727
rect 37191 37449 37207 37727
rect 36897 19727 37207 37449
rect 36897 19449 36913 19727
rect 37191 19449 37207 19727
rect 36897 1727 37207 19449
rect 36897 1449 36913 1727
rect 37191 1449 37207 1727
rect 36897 -173 37207 1449
rect 36897 -451 36913 -173
rect 37191 -451 37207 -173
rect 36897 -947 37207 -451
rect 38757 345587 39067 353101
rect 38757 345309 38773 345587
rect 39051 345309 39067 345587
rect 38757 327587 39067 345309
rect 38757 327309 38773 327587
rect 39051 327309 39067 327587
rect 38757 309587 39067 327309
rect 38757 309309 38773 309587
rect 39051 309309 39067 309587
rect 38757 291587 39067 309309
rect 38757 291309 38773 291587
rect 39051 291309 39067 291587
rect 38757 273587 39067 291309
rect 38757 273309 38773 273587
rect 39051 273309 39067 273587
rect 38757 255587 39067 273309
rect 38757 255309 38773 255587
rect 39051 255309 39067 255587
rect 38757 237587 39067 255309
rect 38757 237309 38773 237587
rect 39051 237309 39067 237587
rect 38757 219587 39067 237309
rect 38757 219309 38773 219587
rect 39051 219309 39067 219587
rect 38757 201587 39067 219309
rect 38757 201309 38773 201587
rect 39051 201309 39067 201587
rect 38757 183587 39067 201309
rect 38757 183309 38773 183587
rect 39051 183309 39067 183587
rect 38757 165587 39067 183309
rect 38757 165309 38773 165587
rect 39051 165309 39067 165587
rect 38757 147587 39067 165309
rect 38757 147309 38773 147587
rect 39051 147309 39067 147587
rect 38757 129587 39067 147309
rect 38757 129309 38773 129587
rect 39051 129309 39067 129587
rect 38757 111587 39067 129309
rect 38757 111309 38773 111587
rect 39051 111309 39067 111587
rect 38757 93587 39067 111309
rect 38757 93309 38773 93587
rect 39051 93309 39067 93587
rect 38757 75587 39067 93309
rect 38757 75309 38773 75587
rect 39051 75309 39067 75587
rect 38757 57587 39067 75309
rect 38757 57309 38773 57587
rect 39051 57309 39067 57587
rect 38757 39587 39067 57309
rect 38757 39309 38773 39587
rect 39051 39309 39067 39587
rect 38757 21587 39067 39309
rect 38757 21309 38773 21587
rect 39051 21309 39067 21587
rect 38757 3587 39067 21309
rect 38757 3309 38773 3587
rect 39051 3309 39067 3587
rect 38757 -1133 39067 3309
rect 38757 -1411 38773 -1133
rect 39051 -1411 39067 -1133
rect 38757 -1907 39067 -1411
rect 40617 347447 40927 354061
rect 40617 347169 40633 347447
rect 40911 347169 40927 347447
rect 40617 329447 40927 347169
rect 40617 329169 40633 329447
rect 40911 329169 40927 329447
rect 40617 311447 40927 329169
rect 40617 311169 40633 311447
rect 40911 311169 40927 311447
rect 40617 293447 40927 311169
rect 40617 293169 40633 293447
rect 40911 293169 40927 293447
rect 40617 275447 40927 293169
rect 40617 275169 40633 275447
rect 40911 275169 40927 275447
rect 40617 257447 40927 275169
rect 40617 257169 40633 257447
rect 40911 257169 40927 257447
rect 40617 239447 40927 257169
rect 40617 239169 40633 239447
rect 40911 239169 40927 239447
rect 40617 221447 40927 239169
rect 40617 221169 40633 221447
rect 40911 221169 40927 221447
rect 40617 203447 40927 221169
rect 40617 203169 40633 203447
rect 40911 203169 40927 203447
rect 40617 185447 40927 203169
rect 40617 185169 40633 185447
rect 40911 185169 40927 185447
rect 40617 167447 40927 185169
rect 40617 167169 40633 167447
rect 40911 167169 40927 167447
rect 40617 149447 40927 167169
rect 40617 149169 40633 149447
rect 40911 149169 40927 149447
rect 40617 131447 40927 149169
rect 40617 131169 40633 131447
rect 40911 131169 40927 131447
rect 40617 113447 40927 131169
rect 40617 113169 40633 113447
rect 40911 113169 40927 113447
rect 40617 95447 40927 113169
rect 40617 95169 40633 95447
rect 40911 95169 40927 95447
rect 40617 77447 40927 95169
rect 40617 77169 40633 77447
rect 40911 77169 40927 77447
rect 40617 59447 40927 77169
rect 40617 59169 40633 59447
rect 40911 59169 40927 59447
rect 40617 41447 40927 59169
rect 40617 41169 40633 41447
rect 40911 41169 40927 41447
rect 40617 23447 40927 41169
rect 40617 23169 40633 23447
rect 40911 23169 40927 23447
rect 40617 5447 40927 23169
rect 40617 5169 40633 5447
rect 40911 5169 40927 5447
rect 40617 -2093 40927 5169
rect 40617 -2371 40633 -2093
rect 40911 -2371 40927 -2093
rect 40617 -2867 40927 -2371
rect 42477 349307 42787 355021
rect 51477 355779 51787 355795
rect 51477 355501 51493 355779
rect 51771 355501 51787 355779
rect 49617 354819 49927 354835
rect 49617 354541 49633 354819
rect 49911 354541 49927 354819
rect 47757 353859 48067 353875
rect 47757 353581 47773 353859
rect 48051 353581 48067 353859
rect 42477 349029 42493 349307
rect 42771 349029 42787 349307
rect 42477 331307 42787 349029
rect 42477 331029 42493 331307
rect 42771 331029 42787 331307
rect 42477 313307 42787 331029
rect 42477 313029 42493 313307
rect 42771 313029 42787 313307
rect 42477 295307 42787 313029
rect 42477 295029 42493 295307
rect 42771 295029 42787 295307
rect 42477 277307 42787 295029
rect 42477 277029 42493 277307
rect 42771 277029 42787 277307
rect 42477 259307 42787 277029
rect 42477 259029 42493 259307
rect 42771 259029 42787 259307
rect 42477 241307 42787 259029
rect 42477 241029 42493 241307
rect 42771 241029 42787 241307
rect 42477 223307 42787 241029
rect 42477 223029 42493 223307
rect 42771 223029 42787 223307
rect 42477 205307 42787 223029
rect 42477 205029 42493 205307
rect 42771 205029 42787 205307
rect 42477 187307 42787 205029
rect 42477 187029 42493 187307
rect 42771 187029 42787 187307
rect 42477 169307 42787 187029
rect 42477 169029 42493 169307
rect 42771 169029 42787 169307
rect 42477 151307 42787 169029
rect 42477 151029 42493 151307
rect 42771 151029 42787 151307
rect 42477 133307 42787 151029
rect 42477 133029 42493 133307
rect 42771 133029 42787 133307
rect 42477 115307 42787 133029
rect 42477 115029 42493 115307
rect 42771 115029 42787 115307
rect 42477 97307 42787 115029
rect 42477 97029 42493 97307
rect 42771 97029 42787 97307
rect 42477 79307 42787 97029
rect 42477 79029 42493 79307
rect 42771 79029 42787 79307
rect 42477 61307 42787 79029
rect 42477 61029 42493 61307
rect 42771 61029 42787 61307
rect 42477 43307 42787 61029
rect 42477 43029 42493 43307
rect 42771 43029 42787 43307
rect 42477 25307 42787 43029
rect 42477 25029 42493 25307
rect 42771 25029 42787 25307
rect 42477 7307 42787 25029
rect 42477 7029 42493 7307
rect 42771 7029 42787 7307
rect 33477 -3811 33493 -3533
rect 33771 -3811 33787 -3533
rect 33477 -3827 33787 -3811
rect 42477 -3053 42787 7029
rect 45897 352899 46207 352915
rect 45897 352621 45913 352899
rect 46191 352621 46207 352899
rect 45897 334727 46207 352621
rect 45897 334449 45913 334727
rect 46191 334449 46207 334727
rect 45897 316727 46207 334449
rect 45897 316449 45913 316727
rect 46191 316449 46207 316727
rect 45897 298727 46207 316449
rect 45897 298449 45913 298727
rect 46191 298449 46207 298727
rect 45897 280727 46207 298449
rect 45897 280449 45913 280727
rect 46191 280449 46207 280727
rect 45897 262727 46207 280449
rect 45897 262449 45913 262727
rect 46191 262449 46207 262727
rect 45897 244727 46207 262449
rect 45897 244449 45913 244727
rect 46191 244449 46207 244727
rect 45897 226727 46207 244449
rect 45897 226449 45913 226727
rect 46191 226449 46207 226727
rect 45897 208727 46207 226449
rect 45897 208449 45913 208727
rect 46191 208449 46207 208727
rect 45897 190727 46207 208449
rect 45897 190449 45913 190727
rect 46191 190449 46207 190727
rect 45897 172727 46207 190449
rect 45897 172449 45913 172727
rect 46191 172449 46207 172727
rect 45897 154727 46207 172449
rect 45897 154449 45913 154727
rect 46191 154449 46207 154727
rect 45897 136727 46207 154449
rect 45897 136449 45913 136727
rect 46191 136449 46207 136727
rect 45897 118727 46207 136449
rect 45897 118449 45913 118727
rect 46191 118449 46207 118727
rect 45897 100727 46207 118449
rect 45897 100449 45913 100727
rect 46191 100449 46207 100727
rect 45897 82727 46207 100449
rect 45897 82449 45913 82727
rect 46191 82449 46207 82727
rect 45897 64727 46207 82449
rect 45897 64449 45913 64727
rect 46191 64449 46207 64727
rect 45897 46727 46207 64449
rect 45897 46449 45913 46727
rect 46191 46449 46207 46727
rect 45897 28727 46207 46449
rect 45897 28449 45913 28727
rect 46191 28449 46207 28727
rect 45897 10727 46207 28449
rect 45897 10449 45913 10727
rect 46191 10449 46207 10727
rect 45897 -653 46207 10449
rect 45897 -931 45913 -653
rect 46191 -931 46207 -653
rect 45897 -947 46207 -931
rect 47757 336587 48067 353581
rect 47757 336309 47773 336587
rect 48051 336309 48067 336587
rect 47757 318587 48067 336309
rect 47757 318309 47773 318587
rect 48051 318309 48067 318587
rect 47757 300587 48067 318309
rect 47757 300309 47773 300587
rect 48051 300309 48067 300587
rect 47757 282587 48067 300309
rect 47757 282309 47773 282587
rect 48051 282309 48067 282587
rect 47757 264587 48067 282309
rect 47757 264309 47773 264587
rect 48051 264309 48067 264587
rect 47757 246587 48067 264309
rect 47757 246309 47773 246587
rect 48051 246309 48067 246587
rect 47757 228587 48067 246309
rect 47757 228309 47773 228587
rect 48051 228309 48067 228587
rect 47757 210587 48067 228309
rect 47757 210309 47773 210587
rect 48051 210309 48067 210587
rect 47757 192587 48067 210309
rect 47757 192309 47773 192587
rect 48051 192309 48067 192587
rect 47757 174587 48067 192309
rect 47757 174309 47773 174587
rect 48051 174309 48067 174587
rect 47757 156587 48067 174309
rect 47757 156309 47773 156587
rect 48051 156309 48067 156587
rect 47757 138587 48067 156309
rect 47757 138309 47773 138587
rect 48051 138309 48067 138587
rect 47757 120587 48067 138309
rect 47757 120309 47773 120587
rect 48051 120309 48067 120587
rect 47757 102587 48067 120309
rect 47757 102309 47773 102587
rect 48051 102309 48067 102587
rect 47757 84587 48067 102309
rect 47757 84309 47773 84587
rect 48051 84309 48067 84587
rect 47757 66587 48067 84309
rect 47757 66309 47773 66587
rect 48051 66309 48067 66587
rect 47757 48587 48067 66309
rect 47757 48309 47773 48587
rect 48051 48309 48067 48587
rect 47757 30587 48067 48309
rect 47757 30309 47773 30587
rect 48051 30309 48067 30587
rect 47757 12587 48067 30309
rect 47757 12309 47773 12587
rect 48051 12309 48067 12587
rect 47757 -1613 48067 12309
rect 47757 -1891 47773 -1613
rect 48051 -1891 48067 -1613
rect 47757 -1907 48067 -1891
rect 49617 338447 49927 354541
rect 49617 338169 49633 338447
rect 49911 338169 49927 338447
rect 49617 320447 49927 338169
rect 49617 320169 49633 320447
rect 49911 320169 49927 320447
rect 49617 302447 49927 320169
rect 49617 302169 49633 302447
rect 49911 302169 49927 302447
rect 49617 284447 49927 302169
rect 49617 284169 49633 284447
rect 49911 284169 49927 284447
rect 49617 266447 49927 284169
rect 49617 266169 49633 266447
rect 49911 266169 49927 266447
rect 49617 248447 49927 266169
rect 49617 248169 49633 248447
rect 49911 248169 49927 248447
rect 49617 230447 49927 248169
rect 49617 230169 49633 230447
rect 49911 230169 49927 230447
rect 49617 212447 49927 230169
rect 49617 212169 49633 212447
rect 49911 212169 49927 212447
rect 49617 194447 49927 212169
rect 49617 194169 49633 194447
rect 49911 194169 49927 194447
rect 49617 176447 49927 194169
rect 49617 176169 49633 176447
rect 49911 176169 49927 176447
rect 49617 158447 49927 176169
rect 49617 158169 49633 158447
rect 49911 158169 49927 158447
rect 49617 140447 49927 158169
rect 49617 140169 49633 140447
rect 49911 140169 49927 140447
rect 49617 122447 49927 140169
rect 49617 122169 49633 122447
rect 49911 122169 49927 122447
rect 49617 104447 49927 122169
rect 49617 104169 49633 104447
rect 49911 104169 49927 104447
rect 49617 86447 49927 104169
rect 49617 86169 49633 86447
rect 49911 86169 49927 86447
rect 49617 68447 49927 86169
rect 49617 68169 49633 68447
rect 49911 68169 49927 68447
rect 49617 50447 49927 68169
rect 49617 50169 49633 50447
rect 49911 50169 49927 50447
rect 49617 32447 49927 50169
rect 49617 32169 49633 32447
rect 49911 32169 49927 32447
rect 49617 14447 49927 32169
rect 49617 14169 49633 14447
rect 49911 14169 49927 14447
rect 49617 -2573 49927 14169
rect 49617 -2851 49633 -2573
rect 49911 -2851 49927 -2573
rect 49617 -2867 49927 -2851
rect 51477 340307 51787 355501
rect 60477 355299 60787 355795
rect 60477 355021 60493 355299
rect 60771 355021 60787 355299
rect 58617 354339 58927 354835
rect 58617 354061 58633 354339
rect 58911 354061 58927 354339
rect 56757 353379 57067 353875
rect 56757 353101 56773 353379
rect 57051 353101 57067 353379
rect 51477 340029 51493 340307
rect 51771 340029 51787 340307
rect 51477 322307 51787 340029
rect 51477 322029 51493 322307
rect 51771 322029 51787 322307
rect 51477 304307 51787 322029
rect 51477 304029 51493 304307
rect 51771 304029 51787 304307
rect 51477 286307 51787 304029
rect 51477 286029 51493 286307
rect 51771 286029 51787 286307
rect 51477 268307 51787 286029
rect 51477 268029 51493 268307
rect 51771 268029 51787 268307
rect 51477 250307 51787 268029
rect 51477 250029 51493 250307
rect 51771 250029 51787 250307
rect 51477 232307 51787 250029
rect 51477 232029 51493 232307
rect 51771 232029 51787 232307
rect 51477 214307 51787 232029
rect 51477 214029 51493 214307
rect 51771 214029 51787 214307
rect 51477 196307 51787 214029
rect 51477 196029 51493 196307
rect 51771 196029 51787 196307
rect 51477 178307 51787 196029
rect 51477 178029 51493 178307
rect 51771 178029 51787 178307
rect 51477 160307 51787 178029
rect 51477 160029 51493 160307
rect 51771 160029 51787 160307
rect 51477 142307 51787 160029
rect 51477 142029 51493 142307
rect 51771 142029 51787 142307
rect 51477 124307 51787 142029
rect 51477 124029 51493 124307
rect 51771 124029 51787 124307
rect 51477 106307 51787 124029
rect 51477 106029 51493 106307
rect 51771 106029 51787 106307
rect 51477 88307 51787 106029
rect 51477 88029 51493 88307
rect 51771 88029 51787 88307
rect 51477 70307 51787 88029
rect 51477 70029 51493 70307
rect 51771 70029 51787 70307
rect 51477 52307 51787 70029
rect 51477 52029 51493 52307
rect 51771 52029 51787 52307
rect 51477 34307 51787 52029
rect 51477 34029 51493 34307
rect 51771 34029 51787 34307
rect 51477 16307 51787 34029
rect 51477 16029 51493 16307
rect 51771 16029 51787 16307
rect 42477 -3331 42493 -3053
rect 42771 -3331 42787 -3053
rect 42477 -3827 42787 -3331
rect 51477 -3533 51787 16029
rect 54897 352419 55207 352915
rect 54897 352141 54913 352419
rect 55191 352141 55207 352419
rect 54897 343727 55207 352141
rect 54897 343449 54913 343727
rect 55191 343449 55207 343727
rect 54897 325727 55207 343449
rect 54897 325449 54913 325727
rect 55191 325449 55207 325727
rect 54897 307727 55207 325449
rect 54897 307449 54913 307727
rect 55191 307449 55207 307727
rect 54897 289727 55207 307449
rect 54897 289449 54913 289727
rect 55191 289449 55207 289727
rect 54897 271727 55207 289449
rect 54897 271449 54913 271727
rect 55191 271449 55207 271727
rect 54897 253727 55207 271449
rect 54897 253449 54913 253727
rect 55191 253449 55207 253727
rect 54897 235727 55207 253449
rect 54897 235449 54913 235727
rect 55191 235449 55207 235727
rect 54897 217727 55207 235449
rect 54897 217449 54913 217727
rect 55191 217449 55207 217727
rect 54897 199727 55207 217449
rect 54897 199449 54913 199727
rect 55191 199449 55207 199727
rect 54897 181727 55207 199449
rect 54897 181449 54913 181727
rect 55191 181449 55207 181727
rect 54897 163727 55207 181449
rect 54897 163449 54913 163727
rect 55191 163449 55207 163727
rect 54897 145727 55207 163449
rect 54897 145449 54913 145727
rect 55191 145449 55207 145727
rect 54897 127727 55207 145449
rect 54897 127449 54913 127727
rect 55191 127449 55207 127727
rect 54897 109727 55207 127449
rect 54897 109449 54913 109727
rect 55191 109449 55207 109727
rect 54897 91727 55207 109449
rect 54897 91449 54913 91727
rect 55191 91449 55207 91727
rect 54897 73727 55207 91449
rect 54897 73449 54913 73727
rect 55191 73449 55207 73727
rect 54897 55727 55207 73449
rect 54897 55449 54913 55727
rect 55191 55449 55207 55727
rect 54897 37727 55207 55449
rect 54897 37449 54913 37727
rect 55191 37449 55207 37727
rect 54897 19727 55207 37449
rect 54897 19449 54913 19727
rect 55191 19449 55207 19727
rect 54897 1727 55207 19449
rect 54897 1449 54913 1727
rect 55191 1449 55207 1727
rect 54897 -173 55207 1449
rect 54897 -451 54913 -173
rect 55191 -451 55207 -173
rect 54897 -947 55207 -451
rect 56757 345587 57067 353101
rect 56757 345309 56773 345587
rect 57051 345309 57067 345587
rect 56757 327587 57067 345309
rect 56757 327309 56773 327587
rect 57051 327309 57067 327587
rect 56757 309587 57067 327309
rect 56757 309309 56773 309587
rect 57051 309309 57067 309587
rect 56757 291587 57067 309309
rect 56757 291309 56773 291587
rect 57051 291309 57067 291587
rect 56757 273587 57067 291309
rect 56757 273309 56773 273587
rect 57051 273309 57067 273587
rect 56757 255587 57067 273309
rect 56757 255309 56773 255587
rect 57051 255309 57067 255587
rect 56757 237587 57067 255309
rect 56757 237309 56773 237587
rect 57051 237309 57067 237587
rect 56757 219587 57067 237309
rect 56757 219309 56773 219587
rect 57051 219309 57067 219587
rect 56757 201587 57067 219309
rect 56757 201309 56773 201587
rect 57051 201309 57067 201587
rect 56757 183587 57067 201309
rect 56757 183309 56773 183587
rect 57051 183309 57067 183587
rect 56757 165587 57067 183309
rect 56757 165309 56773 165587
rect 57051 165309 57067 165587
rect 56757 147587 57067 165309
rect 56757 147309 56773 147587
rect 57051 147309 57067 147587
rect 56757 129587 57067 147309
rect 56757 129309 56773 129587
rect 57051 129309 57067 129587
rect 56757 111587 57067 129309
rect 56757 111309 56773 111587
rect 57051 111309 57067 111587
rect 56757 93587 57067 111309
rect 56757 93309 56773 93587
rect 57051 93309 57067 93587
rect 56757 75587 57067 93309
rect 56757 75309 56773 75587
rect 57051 75309 57067 75587
rect 56757 57587 57067 75309
rect 56757 57309 56773 57587
rect 57051 57309 57067 57587
rect 56757 39587 57067 57309
rect 56757 39309 56773 39587
rect 57051 39309 57067 39587
rect 56757 21587 57067 39309
rect 56757 21309 56773 21587
rect 57051 21309 57067 21587
rect 56757 3587 57067 21309
rect 56757 3309 56773 3587
rect 57051 3309 57067 3587
rect 56757 -1133 57067 3309
rect 56757 -1411 56773 -1133
rect 57051 -1411 57067 -1133
rect 56757 -1907 57067 -1411
rect 58617 347447 58927 354061
rect 58617 347169 58633 347447
rect 58911 347169 58927 347447
rect 58617 329447 58927 347169
rect 58617 329169 58633 329447
rect 58911 329169 58927 329447
rect 58617 311447 58927 329169
rect 58617 311169 58633 311447
rect 58911 311169 58927 311447
rect 58617 293447 58927 311169
rect 58617 293169 58633 293447
rect 58911 293169 58927 293447
rect 58617 275447 58927 293169
rect 58617 275169 58633 275447
rect 58911 275169 58927 275447
rect 58617 257447 58927 275169
rect 58617 257169 58633 257447
rect 58911 257169 58927 257447
rect 58617 239447 58927 257169
rect 58617 239169 58633 239447
rect 58911 239169 58927 239447
rect 58617 221447 58927 239169
rect 58617 221169 58633 221447
rect 58911 221169 58927 221447
rect 58617 203447 58927 221169
rect 58617 203169 58633 203447
rect 58911 203169 58927 203447
rect 58617 185447 58927 203169
rect 58617 185169 58633 185447
rect 58911 185169 58927 185447
rect 58617 167447 58927 185169
rect 58617 167169 58633 167447
rect 58911 167169 58927 167447
rect 58617 149447 58927 167169
rect 58617 149169 58633 149447
rect 58911 149169 58927 149447
rect 58617 131447 58927 149169
rect 58617 131169 58633 131447
rect 58911 131169 58927 131447
rect 58617 113447 58927 131169
rect 58617 113169 58633 113447
rect 58911 113169 58927 113447
rect 58617 95447 58927 113169
rect 58617 95169 58633 95447
rect 58911 95169 58927 95447
rect 58617 77447 58927 95169
rect 58617 77169 58633 77447
rect 58911 77169 58927 77447
rect 58617 59447 58927 77169
rect 58617 59169 58633 59447
rect 58911 59169 58927 59447
rect 58617 41447 58927 59169
rect 58617 41169 58633 41447
rect 58911 41169 58927 41447
rect 58617 23447 58927 41169
rect 58617 23169 58633 23447
rect 58911 23169 58927 23447
rect 58617 5447 58927 23169
rect 58617 5169 58633 5447
rect 58911 5169 58927 5447
rect 58617 -2093 58927 5169
rect 58617 -2371 58633 -2093
rect 58911 -2371 58927 -2093
rect 58617 -2867 58927 -2371
rect 60477 349307 60787 355021
rect 69477 355779 69787 355795
rect 69477 355501 69493 355779
rect 69771 355501 69787 355779
rect 67617 354819 67927 354835
rect 67617 354541 67633 354819
rect 67911 354541 67927 354819
rect 65757 353859 66067 353875
rect 65757 353581 65773 353859
rect 66051 353581 66067 353859
rect 60477 349029 60493 349307
rect 60771 349029 60787 349307
rect 60477 331307 60787 349029
rect 60477 331029 60493 331307
rect 60771 331029 60787 331307
rect 60477 313307 60787 331029
rect 60477 313029 60493 313307
rect 60771 313029 60787 313307
rect 60477 295307 60787 313029
rect 60477 295029 60493 295307
rect 60771 295029 60787 295307
rect 60477 277307 60787 295029
rect 60477 277029 60493 277307
rect 60771 277029 60787 277307
rect 60477 259307 60787 277029
rect 60477 259029 60493 259307
rect 60771 259029 60787 259307
rect 60477 241307 60787 259029
rect 60477 241029 60493 241307
rect 60771 241029 60787 241307
rect 60477 223307 60787 241029
rect 60477 223029 60493 223307
rect 60771 223029 60787 223307
rect 60477 205307 60787 223029
rect 60477 205029 60493 205307
rect 60771 205029 60787 205307
rect 60477 187307 60787 205029
rect 60477 187029 60493 187307
rect 60771 187029 60787 187307
rect 60477 169307 60787 187029
rect 60477 169029 60493 169307
rect 60771 169029 60787 169307
rect 60477 151307 60787 169029
rect 60477 151029 60493 151307
rect 60771 151029 60787 151307
rect 60477 133307 60787 151029
rect 60477 133029 60493 133307
rect 60771 133029 60787 133307
rect 60477 115307 60787 133029
rect 60477 115029 60493 115307
rect 60771 115029 60787 115307
rect 60477 97307 60787 115029
rect 60477 97029 60493 97307
rect 60771 97029 60787 97307
rect 60477 79307 60787 97029
rect 60477 79029 60493 79307
rect 60771 79029 60787 79307
rect 60477 61307 60787 79029
rect 60477 61029 60493 61307
rect 60771 61029 60787 61307
rect 60477 43307 60787 61029
rect 60477 43029 60493 43307
rect 60771 43029 60787 43307
rect 60477 25307 60787 43029
rect 60477 25029 60493 25307
rect 60771 25029 60787 25307
rect 60477 7307 60787 25029
rect 60477 7029 60493 7307
rect 60771 7029 60787 7307
rect 51477 -3811 51493 -3533
rect 51771 -3811 51787 -3533
rect 51477 -3827 51787 -3811
rect 60477 -3053 60787 7029
rect 63897 352899 64207 352915
rect 63897 352621 63913 352899
rect 64191 352621 64207 352899
rect 63897 334727 64207 352621
rect 63897 334449 63913 334727
rect 64191 334449 64207 334727
rect 63897 316727 64207 334449
rect 63897 316449 63913 316727
rect 64191 316449 64207 316727
rect 63897 298727 64207 316449
rect 63897 298449 63913 298727
rect 64191 298449 64207 298727
rect 63897 280727 64207 298449
rect 63897 280449 63913 280727
rect 64191 280449 64207 280727
rect 63897 262727 64207 280449
rect 63897 262449 63913 262727
rect 64191 262449 64207 262727
rect 63897 244727 64207 262449
rect 63897 244449 63913 244727
rect 64191 244449 64207 244727
rect 63897 226727 64207 244449
rect 63897 226449 63913 226727
rect 64191 226449 64207 226727
rect 63897 208727 64207 226449
rect 63897 208449 63913 208727
rect 64191 208449 64207 208727
rect 63897 190727 64207 208449
rect 63897 190449 63913 190727
rect 64191 190449 64207 190727
rect 63897 172727 64207 190449
rect 63897 172449 63913 172727
rect 64191 172449 64207 172727
rect 63897 154727 64207 172449
rect 63897 154449 63913 154727
rect 64191 154449 64207 154727
rect 63897 136727 64207 154449
rect 63897 136449 63913 136727
rect 64191 136449 64207 136727
rect 63897 118727 64207 136449
rect 63897 118449 63913 118727
rect 64191 118449 64207 118727
rect 63897 100727 64207 118449
rect 63897 100449 63913 100727
rect 64191 100449 64207 100727
rect 63897 82727 64207 100449
rect 63897 82449 63913 82727
rect 64191 82449 64207 82727
rect 63897 64727 64207 82449
rect 63897 64449 63913 64727
rect 64191 64449 64207 64727
rect 63897 46727 64207 64449
rect 63897 46449 63913 46727
rect 64191 46449 64207 46727
rect 63897 28727 64207 46449
rect 63897 28449 63913 28727
rect 64191 28449 64207 28727
rect 63897 10727 64207 28449
rect 63897 10449 63913 10727
rect 64191 10449 64207 10727
rect 63897 -653 64207 10449
rect 63897 -931 63913 -653
rect 64191 -931 64207 -653
rect 63897 -947 64207 -931
rect 65757 336587 66067 353581
rect 65757 336309 65773 336587
rect 66051 336309 66067 336587
rect 65757 318587 66067 336309
rect 65757 318309 65773 318587
rect 66051 318309 66067 318587
rect 65757 300587 66067 318309
rect 65757 300309 65773 300587
rect 66051 300309 66067 300587
rect 65757 282587 66067 300309
rect 65757 282309 65773 282587
rect 66051 282309 66067 282587
rect 65757 264587 66067 282309
rect 65757 264309 65773 264587
rect 66051 264309 66067 264587
rect 65757 246587 66067 264309
rect 65757 246309 65773 246587
rect 66051 246309 66067 246587
rect 65757 228587 66067 246309
rect 65757 228309 65773 228587
rect 66051 228309 66067 228587
rect 65757 210587 66067 228309
rect 65757 210309 65773 210587
rect 66051 210309 66067 210587
rect 65757 192587 66067 210309
rect 65757 192309 65773 192587
rect 66051 192309 66067 192587
rect 65757 174587 66067 192309
rect 65757 174309 65773 174587
rect 66051 174309 66067 174587
rect 65757 156587 66067 174309
rect 65757 156309 65773 156587
rect 66051 156309 66067 156587
rect 65757 138587 66067 156309
rect 65757 138309 65773 138587
rect 66051 138309 66067 138587
rect 65757 120587 66067 138309
rect 65757 120309 65773 120587
rect 66051 120309 66067 120587
rect 65757 102587 66067 120309
rect 65757 102309 65773 102587
rect 66051 102309 66067 102587
rect 65757 84587 66067 102309
rect 65757 84309 65773 84587
rect 66051 84309 66067 84587
rect 65757 66587 66067 84309
rect 65757 66309 65773 66587
rect 66051 66309 66067 66587
rect 65757 48587 66067 66309
rect 65757 48309 65773 48587
rect 66051 48309 66067 48587
rect 65757 30587 66067 48309
rect 65757 30309 65773 30587
rect 66051 30309 66067 30587
rect 65757 12587 66067 30309
rect 65757 12309 65773 12587
rect 66051 12309 66067 12587
rect 65757 -1613 66067 12309
rect 65757 -1891 65773 -1613
rect 66051 -1891 66067 -1613
rect 65757 -1907 66067 -1891
rect 67617 338447 67927 354541
rect 67617 338169 67633 338447
rect 67911 338169 67927 338447
rect 67617 320447 67927 338169
rect 67617 320169 67633 320447
rect 67911 320169 67927 320447
rect 67617 302447 67927 320169
rect 67617 302169 67633 302447
rect 67911 302169 67927 302447
rect 67617 284447 67927 302169
rect 67617 284169 67633 284447
rect 67911 284169 67927 284447
rect 67617 266447 67927 284169
rect 67617 266169 67633 266447
rect 67911 266169 67927 266447
rect 67617 248447 67927 266169
rect 67617 248169 67633 248447
rect 67911 248169 67927 248447
rect 67617 230447 67927 248169
rect 67617 230169 67633 230447
rect 67911 230169 67927 230447
rect 67617 212447 67927 230169
rect 67617 212169 67633 212447
rect 67911 212169 67927 212447
rect 67617 194447 67927 212169
rect 67617 194169 67633 194447
rect 67911 194169 67927 194447
rect 67617 176447 67927 194169
rect 67617 176169 67633 176447
rect 67911 176169 67927 176447
rect 67617 158447 67927 176169
rect 67617 158169 67633 158447
rect 67911 158169 67927 158447
rect 67617 140447 67927 158169
rect 67617 140169 67633 140447
rect 67911 140169 67927 140447
rect 67617 122447 67927 140169
rect 67617 122169 67633 122447
rect 67911 122169 67927 122447
rect 67617 104447 67927 122169
rect 67617 104169 67633 104447
rect 67911 104169 67927 104447
rect 67617 86447 67927 104169
rect 67617 86169 67633 86447
rect 67911 86169 67927 86447
rect 67617 68447 67927 86169
rect 67617 68169 67633 68447
rect 67911 68169 67927 68447
rect 67617 50447 67927 68169
rect 67617 50169 67633 50447
rect 67911 50169 67927 50447
rect 67617 32447 67927 50169
rect 67617 32169 67633 32447
rect 67911 32169 67927 32447
rect 67617 14447 67927 32169
rect 67617 14169 67633 14447
rect 67911 14169 67927 14447
rect 67617 -2573 67927 14169
rect 67617 -2851 67633 -2573
rect 67911 -2851 67927 -2573
rect 67617 -2867 67927 -2851
rect 69477 340307 69787 355501
rect 78477 355299 78787 355795
rect 78477 355021 78493 355299
rect 78771 355021 78787 355299
rect 76617 354339 76927 354835
rect 76617 354061 76633 354339
rect 76911 354061 76927 354339
rect 74757 353379 75067 353875
rect 74757 353101 74773 353379
rect 75051 353101 75067 353379
rect 69477 340029 69493 340307
rect 69771 340029 69787 340307
rect 69477 322307 69787 340029
rect 69477 322029 69493 322307
rect 69771 322029 69787 322307
rect 69477 304307 69787 322029
rect 69477 304029 69493 304307
rect 69771 304029 69787 304307
rect 69477 286307 69787 304029
rect 69477 286029 69493 286307
rect 69771 286029 69787 286307
rect 69477 268307 69787 286029
rect 69477 268029 69493 268307
rect 69771 268029 69787 268307
rect 69477 250307 69787 268029
rect 69477 250029 69493 250307
rect 69771 250029 69787 250307
rect 69477 232307 69787 250029
rect 69477 232029 69493 232307
rect 69771 232029 69787 232307
rect 69477 214307 69787 232029
rect 69477 214029 69493 214307
rect 69771 214029 69787 214307
rect 69477 196307 69787 214029
rect 69477 196029 69493 196307
rect 69771 196029 69787 196307
rect 69477 178307 69787 196029
rect 69477 178029 69493 178307
rect 69771 178029 69787 178307
rect 69477 160307 69787 178029
rect 69477 160029 69493 160307
rect 69771 160029 69787 160307
rect 69477 142307 69787 160029
rect 69477 142029 69493 142307
rect 69771 142029 69787 142307
rect 69477 124307 69787 142029
rect 69477 124029 69493 124307
rect 69771 124029 69787 124307
rect 69477 106307 69787 124029
rect 69477 106029 69493 106307
rect 69771 106029 69787 106307
rect 69477 88307 69787 106029
rect 69477 88029 69493 88307
rect 69771 88029 69787 88307
rect 69477 70307 69787 88029
rect 69477 70029 69493 70307
rect 69771 70029 69787 70307
rect 69477 52307 69787 70029
rect 69477 52029 69493 52307
rect 69771 52029 69787 52307
rect 69477 34307 69787 52029
rect 69477 34029 69493 34307
rect 69771 34029 69787 34307
rect 69477 16307 69787 34029
rect 69477 16029 69493 16307
rect 69771 16029 69787 16307
rect 60477 -3331 60493 -3053
rect 60771 -3331 60787 -3053
rect 60477 -3827 60787 -3331
rect 69477 -3533 69787 16029
rect 72897 352419 73207 352915
rect 72897 352141 72913 352419
rect 73191 352141 73207 352419
rect 72897 343727 73207 352141
rect 72897 343449 72913 343727
rect 73191 343449 73207 343727
rect 72897 325727 73207 343449
rect 72897 325449 72913 325727
rect 73191 325449 73207 325727
rect 72897 307727 73207 325449
rect 72897 307449 72913 307727
rect 73191 307449 73207 307727
rect 72897 289727 73207 307449
rect 72897 289449 72913 289727
rect 73191 289449 73207 289727
rect 72897 271727 73207 289449
rect 72897 271449 72913 271727
rect 73191 271449 73207 271727
rect 72897 253727 73207 271449
rect 72897 253449 72913 253727
rect 73191 253449 73207 253727
rect 72897 235727 73207 253449
rect 72897 235449 72913 235727
rect 73191 235449 73207 235727
rect 72897 217727 73207 235449
rect 72897 217449 72913 217727
rect 73191 217449 73207 217727
rect 72897 199727 73207 217449
rect 72897 199449 72913 199727
rect 73191 199449 73207 199727
rect 72897 181727 73207 199449
rect 72897 181449 72913 181727
rect 73191 181449 73207 181727
rect 72897 163727 73207 181449
rect 72897 163449 72913 163727
rect 73191 163449 73207 163727
rect 72897 145727 73207 163449
rect 72897 145449 72913 145727
rect 73191 145449 73207 145727
rect 72897 127727 73207 145449
rect 72897 127449 72913 127727
rect 73191 127449 73207 127727
rect 72897 109727 73207 127449
rect 72897 109449 72913 109727
rect 73191 109449 73207 109727
rect 72897 91727 73207 109449
rect 72897 91449 72913 91727
rect 73191 91449 73207 91727
rect 72897 73727 73207 91449
rect 72897 73449 72913 73727
rect 73191 73449 73207 73727
rect 72897 55727 73207 73449
rect 72897 55449 72913 55727
rect 73191 55449 73207 55727
rect 72897 37727 73207 55449
rect 72897 37449 72913 37727
rect 73191 37449 73207 37727
rect 72897 19727 73207 37449
rect 72897 19449 72913 19727
rect 73191 19449 73207 19727
rect 72897 1727 73207 19449
rect 72897 1449 72913 1727
rect 73191 1449 73207 1727
rect 72897 -173 73207 1449
rect 72897 -451 72913 -173
rect 73191 -451 73207 -173
rect 72897 -947 73207 -451
rect 74757 345587 75067 353101
rect 74757 345309 74773 345587
rect 75051 345309 75067 345587
rect 74757 327587 75067 345309
rect 74757 327309 74773 327587
rect 75051 327309 75067 327587
rect 74757 309587 75067 327309
rect 74757 309309 74773 309587
rect 75051 309309 75067 309587
rect 74757 291587 75067 309309
rect 74757 291309 74773 291587
rect 75051 291309 75067 291587
rect 74757 273587 75067 291309
rect 74757 273309 74773 273587
rect 75051 273309 75067 273587
rect 74757 255587 75067 273309
rect 74757 255309 74773 255587
rect 75051 255309 75067 255587
rect 74757 237587 75067 255309
rect 74757 237309 74773 237587
rect 75051 237309 75067 237587
rect 74757 219587 75067 237309
rect 74757 219309 74773 219587
rect 75051 219309 75067 219587
rect 74757 201587 75067 219309
rect 74757 201309 74773 201587
rect 75051 201309 75067 201587
rect 74757 183587 75067 201309
rect 74757 183309 74773 183587
rect 75051 183309 75067 183587
rect 74757 165587 75067 183309
rect 74757 165309 74773 165587
rect 75051 165309 75067 165587
rect 74757 147587 75067 165309
rect 74757 147309 74773 147587
rect 75051 147309 75067 147587
rect 74757 129587 75067 147309
rect 74757 129309 74773 129587
rect 75051 129309 75067 129587
rect 74757 111587 75067 129309
rect 74757 111309 74773 111587
rect 75051 111309 75067 111587
rect 74757 93587 75067 111309
rect 74757 93309 74773 93587
rect 75051 93309 75067 93587
rect 74757 75587 75067 93309
rect 74757 75309 74773 75587
rect 75051 75309 75067 75587
rect 74757 57587 75067 75309
rect 74757 57309 74773 57587
rect 75051 57309 75067 57587
rect 74757 39587 75067 57309
rect 74757 39309 74773 39587
rect 75051 39309 75067 39587
rect 74757 21587 75067 39309
rect 74757 21309 74773 21587
rect 75051 21309 75067 21587
rect 74757 3587 75067 21309
rect 74757 3309 74773 3587
rect 75051 3309 75067 3587
rect 74757 -1133 75067 3309
rect 74757 -1411 74773 -1133
rect 75051 -1411 75067 -1133
rect 74757 -1907 75067 -1411
rect 76617 347447 76927 354061
rect 76617 347169 76633 347447
rect 76911 347169 76927 347447
rect 76617 329447 76927 347169
rect 76617 329169 76633 329447
rect 76911 329169 76927 329447
rect 76617 311447 76927 329169
rect 76617 311169 76633 311447
rect 76911 311169 76927 311447
rect 76617 293447 76927 311169
rect 76617 293169 76633 293447
rect 76911 293169 76927 293447
rect 76617 275447 76927 293169
rect 76617 275169 76633 275447
rect 76911 275169 76927 275447
rect 76617 257447 76927 275169
rect 76617 257169 76633 257447
rect 76911 257169 76927 257447
rect 76617 239447 76927 257169
rect 76617 239169 76633 239447
rect 76911 239169 76927 239447
rect 76617 221447 76927 239169
rect 76617 221169 76633 221447
rect 76911 221169 76927 221447
rect 76617 203447 76927 221169
rect 76617 203169 76633 203447
rect 76911 203169 76927 203447
rect 76617 185447 76927 203169
rect 76617 185169 76633 185447
rect 76911 185169 76927 185447
rect 76617 167447 76927 185169
rect 76617 167169 76633 167447
rect 76911 167169 76927 167447
rect 76617 149447 76927 167169
rect 76617 149169 76633 149447
rect 76911 149169 76927 149447
rect 76617 131447 76927 149169
rect 76617 131169 76633 131447
rect 76911 131169 76927 131447
rect 76617 113447 76927 131169
rect 76617 113169 76633 113447
rect 76911 113169 76927 113447
rect 76617 95447 76927 113169
rect 76617 95169 76633 95447
rect 76911 95169 76927 95447
rect 76617 77447 76927 95169
rect 76617 77169 76633 77447
rect 76911 77169 76927 77447
rect 76617 59447 76927 77169
rect 76617 59169 76633 59447
rect 76911 59169 76927 59447
rect 76617 41447 76927 59169
rect 76617 41169 76633 41447
rect 76911 41169 76927 41447
rect 76617 23447 76927 41169
rect 76617 23169 76633 23447
rect 76911 23169 76927 23447
rect 76617 5447 76927 23169
rect 76617 5169 76633 5447
rect 76911 5169 76927 5447
rect 76617 -2093 76927 5169
rect 76617 -2371 76633 -2093
rect 76911 -2371 76927 -2093
rect 76617 -2867 76927 -2371
rect 78477 349307 78787 355021
rect 87477 355779 87787 355795
rect 87477 355501 87493 355779
rect 87771 355501 87787 355779
rect 85617 354819 85927 354835
rect 85617 354541 85633 354819
rect 85911 354541 85927 354819
rect 83757 353859 84067 353875
rect 83757 353581 83773 353859
rect 84051 353581 84067 353859
rect 78477 349029 78493 349307
rect 78771 349029 78787 349307
rect 78477 331307 78787 349029
rect 78477 331029 78493 331307
rect 78771 331029 78787 331307
rect 78477 313307 78787 331029
rect 78477 313029 78493 313307
rect 78771 313029 78787 313307
rect 78477 295307 78787 313029
rect 78477 295029 78493 295307
rect 78771 295029 78787 295307
rect 78477 277307 78787 295029
rect 78477 277029 78493 277307
rect 78771 277029 78787 277307
rect 78477 259307 78787 277029
rect 78477 259029 78493 259307
rect 78771 259029 78787 259307
rect 78477 241307 78787 259029
rect 78477 241029 78493 241307
rect 78771 241029 78787 241307
rect 78477 223307 78787 241029
rect 78477 223029 78493 223307
rect 78771 223029 78787 223307
rect 78477 205307 78787 223029
rect 78477 205029 78493 205307
rect 78771 205029 78787 205307
rect 78477 187307 78787 205029
rect 78477 187029 78493 187307
rect 78771 187029 78787 187307
rect 78477 169307 78787 187029
rect 78477 169029 78493 169307
rect 78771 169029 78787 169307
rect 78477 151307 78787 169029
rect 78477 151029 78493 151307
rect 78771 151029 78787 151307
rect 78477 133307 78787 151029
rect 78477 133029 78493 133307
rect 78771 133029 78787 133307
rect 78477 115307 78787 133029
rect 78477 115029 78493 115307
rect 78771 115029 78787 115307
rect 78477 97307 78787 115029
rect 78477 97029 78493 97307
rect 78771 97029 78787 97307
rect 78477 79307 78787 97029
rect 78477 79029 78493 79307
rect 78771 79029 78787 79307
rect 78477 61307 78787 79029
rect 78477 61029 78493 61307
rect 78771 61029 78787 61307
rect 78477 43307 78787 61029
rect 78477 43029 78493 43307
rect 78771 43029 78787 43307
rect 78477 25307 78787 43029
rect 78477 25029 78493 25307
rect 78771 25029 78787 25307
rect 78477 7307 78787 25029
rect 78477 7029 78493 7307
rect 78771 7029 78787 7307
rect 69477 -3811 69493 -3533
rect 69771 -3811 69787 -3533
rect 69477 -3827 69787 -3811
rect 78477 -3053 78787 7029
rect 81897 352899 82207 352915
rect 81897 352621 81913 352899
rect 82191 352621 82207 352899
rect 81897 334727 82207 352621
rect 81897 334449 81913 334727
rect 82191 334449 82207 334727
rect 81897 316727 82207 334449
rect 81897 316449 81913 316727
rect 82191 316449 82207 316727
rect 81897 298727 82207 316449
rect 81897 298449 81913 298727
rect 82191 298449 82207 298727
rect 81897 280727 82207 298449
rect 81897 280449 81913 280727
rect 82191 280449 82207 280727
rect 81897 262727 82207 280449
rect 81897 262449 81913 262727
rect 82191 262449 82207 262727
rect 81897 244727 82207 262449
rect 81897 244449 81913 244727
rect 82191 244449 82207 244727
rect 81897 226727 82207 244449
rect 81897 226449 81913 226727
rect 82191 226449 82207 226727
rect 81897 208727 82207 226449
rect 81897 208449 81913 208727
rect 82191 208449 82207 208727
rect 81897 190727 82207 208449
rect 81897 190449 81913 190727
rect 82191 190449 82207 190727
rect 81897 172727 82207 190449
rect 81897 172449 81913 172727
rect 82191 172449 82207 172727
rect 81897 154727 82207 172449
rect 81897 154449 81913 154727
rect 82191 154449 82207 154727
rect 81897 136727 82207 154449
rect 81897 136449 81913 136727
rect 82191 136449 82207 136727
rect 81897 118727 82207 136449
rect 81897 118449 81913 118727
rect 82191 118449 82207 118727
rect 81897 100727 82207 118449
rect 81897 100449 81913 100727
rect 82191 100449 82207 100727
rect 81897 82727 82207 100449
rect 81897 82449 81913 82727
rect 82191 82449 82207 82727
rect 81897 64727 82207 82449
rect 81897 64449 81913 64727
rect 82191 64449 82207 64727
rect 81897 46727 82207 64449
rect 81897 46449 81913 46727
rect 82191 46449 82207 46727
rect 81897 28727 82207 46449
rect 81897 28449 81913 28727
rect 82191 28449 82207 28727
rect 81897 10727 82207 28449
rect 81897 10449 81913 10727
rect 82191 10449 82207 10727
rect 81897 -653 82207 10449
rect 81897 -931 81913 -653
rect 82191 -931 82207 -653
rect 81897 -947 82207 -931
rect 83757 336587 84067 353581
rect 83757 336309 83773 336587
rect 84051 336309 84067 336587
rect 83757 318587 84067 336309
rect 83757 318309 83773 318587
rect 84051 318309 84067 318587
rect 83757 300587 84067 318309
rect 83757 300309 83773 300587
rect 84051 300309 84067 300587
rect 83757 282587 84067 300309
rect 83757 282309 83773 282587
rect 84051 282309 84067 282587
rect 83757 264587 84067 282309
rect 83757 264309 83773 264587
rect 84051 264309 84067 264587
rect 83757 246587 84067 264309
rect 83757 246309 83773 246587
rect 84051 246309 84067 246587
rect 83757 228587 84067 246309
rect 83757 228309 83773 228587
rect 84051 228309 84067 228587
rect 83757 210587 84067 228309
rect 83757 210309 83773 210587
rect 84051 210309 84067 210587
rect 83757 192587 84067 210309
rect 83757 192309 83773 192587
rect 84051 192309 84067 192587
rect 83757 174587 84067 192309
rect 83757 174309 83773 174587
rect 84051 174309 84067 174587
rect 83757 156587 84067 174309
rect 83757 156309 83773 156587
rect 84051 156309 84067 156587
rect 83757 138587 84067 156309
rect 83757 138309 83773 138587
rect 84051 138309 84067 138587
rect 83757 120587 84067 138309
rect 83757 120309 83773 120587
rect 84051 120309 84067 120587
rect 83757 102587 84067 120309
rect 83757 102309 83773 102587
rect 84051 102309 84067 102587
rect 83757 84587 84067 102309
rect 83757 84309 83773 84587
rect 84051 84309 84067 84587
rect 83757 66587 84067 84309
rect 83757 66309 83773 66587
rect 84051 66309 84067 66587
rect 83757 48587 84067 66309
rect 83757 48309 83773 48587
rect 84051 48309 84067 48587
rect 83757 30587 84067 48309
rect 83757 30309 83773 30587
rect 84051 30309 84067 30587
rect 83757 12587 84067 30309
rect 83757 12309 83773 12587
rect 84051 12309 84067 12587
rect 83757 -1613 84067 12309
rect 83757 -1891 83773 -1613
rect 84051 -1891 84067 -1613
rect 83757 -1907 84067 -1891
rect 85617 338447 85927 354541
rect 85617 338169 85633 338447
rect 85911 338169 85927 338447
rect 85617 320447 85927 338169
rect 85617 320169 85633 320447
rect 85911 320169 85927 320447
rect 85617 302447 85927 320169
rect 85617 302169 85633 302447
rect 85911 302169 85927 302447
rect 85617 284447 85927 302169
rect 85617 284169 85633 284447
rect 85911 284169 85927 284447
rect 85617 266447 85927 284169
rect 85617 266169 85633 266447
rect 85911 266169 85927 266447
rect 85617 248447 85927 266169
rect 85617 248169 85633 248447
rect 85911 248169 85927 248447
rect 85617 230447 85927 248169
rect 85617 230169 85633 230447
rect 85911 230169 85927 230447
rect 85617 212447 85927 230169
rect 85617 212169 85633 212447
rect 85911 212169 85927 212447
rect 85617 194447 85927 212169
rect 85617 194169 85633 194447
rect 85911 194169 85927 194447
rect 85617 176447 85927 194169
rect 85617 176169 85633 176447
rect 85911 176169 85927 176447
rect 85617 158447 85927 176169
rect 85617 158169 85633 158447
rect 85911 158169 85927 158447
rect 85617 140447 85927 158169
rect 85617 140169 85633 140447
rect 85911 140169 85927 140447
rect 85617 122447 85927 140169
rect 85617 122169 85633 122447
rect 85911 122169 85927 122447
rect 85617 104447 85927 122169
rect 85617 104169 85633 104447
rect 85911 104169 85927 104447
rect 85617 86447 85927 104169
rect 85617 86169 85633 86447
rect 85911 86169 85927 86447
rect 85617 68447 85927 86169
rect 85617 68169 85633 68447
rect 85911 68169 85927 68447
rect 85617 50447 85927 68169
rect 85617 50169 85633 50447
rect 85911 50169 85927 50447
rect 85617 32447 85927 50169
rect 85617 32169 85633 32447
rect 85911 32169 85927 32447
rect 85617 14447 85927 32169
rect 85617 14169 85633 14447
rect 85911 14169 85927 14447
rect 85617 -2573 85927 14169
rect 85617 -2851 85633 -2573
rect 85911 -2851 85927 -2573
rect 85617 -2867 85927 -2851
rect 87477 340307 87787 355501
rect 96477 355299 96787 355795
rect 96477 355021 96493 355299
rect 96771 355021 96787 355299
rect 94617 354339 94927 354835
rect 94617 354061 94633 354339
rect 94911 354061 94927 354339
rect 92757 353379 93067 353875
rect 92757 353101 92773 353379
rect 93051 353101 93067 353379
rect 87477 340029 87493 340307
rect 87771 340029 87787 340307
rect 87477 322307 87787 340029
rect 87477 322029 87493 322307
rect 87771 322029 87787 322307
rect 87477 304307 87787 322029
rect 87477 304029 87493 304307
rect 87771 304029 87787 304307
rect 87477 286307 87787 304029
rect 87477 286029 87493 286307
rect 87771 286029 87787 286307
rect 87477 268307 87787 286029
rect 87477 268029 87493 268307
rect 87771 268029 87787 268307
rect 87477 250307 87787 268029
rect 87477 250029 87493 250307
rect 87771 250029 87787 250307
rect 87477 232307 87787 250029
rect 87477 232029 87493 232307
rect 87771 232029 87787 232307
rect 87477 214307 87787 232029
rect 87477 214029 87493 214307
rect 87771 214029 87787 214307
rect 87477 196307 87787 214029
rect 87477 196029 87493 196307
rect 87771 196029 87787 196307
rect 87477 178307 87787 196029
rect 87477 178029 87493 178307
rect 87771 178029 87787 178307
rect 87477 160307 87787 178029
rect 87477 160029 87493 160307
rect 87771 160029 87787 160307
rect 87477 142307 87787 160029
rect 87477 142029 87493 142307
rect 87771 142029 87787 142307
rect 87477 124307 87787 142029
rect 87477 124029 87493 124307
rect 87771 124029 87787 124307
rect 87477 106307 87787 124029
rect 87477 106029 87493 106307
rect 87771 106029 87787 106307
rect 87477 88307 87787 106029
rect 87477 88029 87493 88307
rect 87771 88029 87787 88307
rect 87477 70307 87787 88029
rect 87477 70029 87493 70307
rect 87771 70029 87787 70307
rect 87477 52307 87787 70029
rect 87477 52029 87493 52307
rect 87771 52029 87787 52307
rect 87477 34307 87787 52029
rect 87477 34029 87493 34307
rect 87771 34029 87787 34307
rect 87477 16307 87787 34029
rect 87477 16029 87493 16307
rect 87771 16029 87787 16307
rect 78477 -3331 78493 -3053
rect 78771 -3331 78787 -3053
rect 78477 -3827 78787 -3331
rect 87477 -3533 87787 16029
rect 90897 352419 91207 352915
rect 90897 352141 90913 352419
rect 91191 352141 91207 352419
rect 90897 343727 91207 352141
rect 90897 343449 90913 343727
rect 91191 343449 91207 343727
rect 90897 325727 91207 343449
rect 90897 325449 90913 325727
rect 91191 325449 91207 325727
rect 90897 307727 91207 325449
rect 90897 307449 90913 307727
rect 91191 307449 91207 307727
rect 90897 289727 91207 307449
rect 90897 289449 90913 289727
rect 91191 289449 91207 289727
rect 90897 271727 91207 289449
rect 90897 271449 90913 271727
rect 91191 271449 91207 271727
rect 90897 253727 91207 271449
rect 90897 253449 90913 253727
rect 91191 253449 91207 253727
rect 90897 235727 91207 253449
rect 90897 235449 90913 235727
rect 91191 235449 91207 235727
rect 90897 217727 91207 235449
rect 90897 217449 90913 217727
rect 91191 217449 91207 217727
rect 90897 199727 91207 217449
rect 90897 199449 90913 199727
rect 91191 199449 91207 199727
rect 90897 181727 91207 199449
rect 90897 181449 90913 181727
rect 91191 181449 91207 181727
rect 90897 163727 91207 181449
rect 90897 163449 90913 163727
rect 91191 163449 91207 163727
rect 90897 145727 91207 163449
rect 90897 145449 90913 145727
rect 91191 145449 91207 145727
rect 90897 127727 91207 145449
rect 90897 127449 90913 127727
rect 91191 127449 91207 127727
rect 90897 109727 91207 127449
rect 90897 109449 90913 109727
rect 91191 109449 91207 109727
rect 90897 91727 91207 109449
rect 90897 91449 90913 91727
rect 91191 91449 91207 91727
rect 90897 73727 91207 91449
rect 90897 73449 90913 73727
rect 91191 73449 91207 73727
rect 90897 55727 91207 73449
rect 90897 55449 90913 55727
rect 91191 55449 91207 55727
rect 90897 37727 91207 55449
rect 90897 37449 90913 37727
rect 91191 37449 91207 37727
rect 90897 19727 91207 37449
rect 90897 19449 90913 19727
rect 91191 19449 91207 19727
rect 90897 1727 91207 19449
rect 90897 1449 90913 1727
rect 91191 1449 91207 1727
rect 90897 -173 91207 1449
rect 90897 -451 90913 -173
rect 91191 -451 91207 -173
rect 90897 -947 91207 -451
rect 92757 345587 93067 353101
rect 92757 345309 92773 345587
rect 93051 345309 93067 345587
rect 92757 327587 93067 345309
rect 92757 327309 92773 327587
rect 93051 327309 93067 327587
rect 92757 309587 93067 327309
rect 92757 309309 92773 309587
rect 93051 309309 93067 309587
rect 92757 291587 93067 309309
rect 92757 291309 92773 291587
rect 93051 291309 93067 291587
rect 92757 273587 93067 291309
rect 92757 273309 92773 273587
rect 93051 273309 93067 273587
rect 92757 255587 93067 273309
rect 92757 255309 92773 255587
rect 93051 255309 93067 255587
rect 92757 237587 93067 255309
rect 92757 237309 92773 237587
rect 93051 237309 93067 237587
rect 92757 219587 93067 237309
rect 92757 219309 92773 219587
rect 93051 219309 93067 219587
rect 92757 201587 93067 219309
rect 92757 201309 92773 201587
rect 93051 201309 93067 201587
rect 92757 183587 93067 201309
rect 92757 183309 92773 183587
rect 93051 183309 93067 183587
rect 92757 165587 93067 183309
rect 92757 165309 92773 165587
rect 93051 165309 93067 165587
rect 92757 147587 93067 165309
rect 92757 147309 92773 147587
rect 93051 147309 93067 147587
rect 92757 129587 93067 147309
rect 92757 129309 92773 129587
rect 93051 129309 93067 129587
rect 92757 111587 93067 129309
rect 92757 111309 92773 111587
rect 93051 111309 93067 111587
rect 92757 93587 93067 111309
rect 92757 93309 92773 93587
rect 93051 93309 93067 93587
rect 92757 75587 93067 93309
rect 92757 75309 92773 75587
rect 93051 75309 93067 75587
rect 92757 57587 93067 75309
rect 92757 57309 92773 57587
rect 93051 57309 93067 57587
rect 92757 39587 93067 57309
rect 92757 39309 92773 39587
rect 93051 39309 93067 39587
rect 92757 21587 93067 39309
rect 92757 21309 92773 21587
rect 93051 21309 93067 21587
rect 92757 3587 93067 21309
rect 92757 3309 92773 3587
rect 93051 3309 93067 3587
rect 92757 -1133 93067 3309
rect 92757 -1411 92773 -1133
rect 93051 -1411 93067 -1133
rect 92757 -1907 93067 -1411
rect 94617 347447 94927 354061
rect 94617 347169 94633 347447
rect 94911 347169 94927 347447
rect 94617 329447 94927 347169
rect 94617 329169 94633 329447
rect 94911 329169 94927 329447
rect 94617 311447 94927 329169
rect 94617 311169 94633 311447
rect 94911 311169 94927 311447
rect 94617 293447 94927 311169
rect 94617 293169 94633 293447
rect 94911 293169 94927 293447
rect 94617 275447 94927 293169
rect 94617 275169 94633 275447
rect 94911 275169 94927 275447
rect 94617 257447 94927 275169
rect 94617 257169 94633 257447
rect 94911 257169 94927 257447
rect 94617 239447 94927 257169
rect 94617 239169 94633 239447
rect 94911 239169 94927 239447
rect 94617 221447 94927 239169
rect 94617 221169 94633 221447
rect 94911 221169 94927 221447
rect 94617 203447 94927 221169
rect 94617 203169 94633 203447
rect 94911 203169 94927 203447
rect 94617 185447 94927 203169
rect 94617 185169 94633 185447
rect 94911 185169 94927 185447
rect 94617 167447 94927 185169
rect 94617 167169 94633 167447
rect 94911 167169 94927 167447
rect 94617 149447 94927 167169
rect 94617 149169 94633 149447
rect 94911 149169 94927 149447
rect 94617 131447 94927 149169
rect 94617 131169 94633 131447
rect 94911 131169 94927 131447
rect 94617 113447 94927 131169
rect 94617 113169 94633 113447
rect 94911 113169 94927 113447
rect 94617 95447 94927 113169
rect 94617 95169 94633 95447
rect 94911 95169 94927 95447
rect 94617 77447 94927 95169
rect 94617 77169 94633 77447
rect 94911 77169 94927 77447
rect 94617 59447 94927 77169
rect 94617 59169 94633 59447
rect 94911 59169 94927 59447
rect 94617 41447 94927 59169
rect 94617 41169 94633 41447
rect 94911 41169 94927 41447
rect 94617 23447 94927 41169
rect 94617 23169 94633 23447
rect 94911 23169 94927 23447
rect 94617 5447 94927 23169
rect 94617 5169 94633 5447
rect 94911 5169 94927 5447
rect 94617 -2093 94927 5169
rect 94617 -2371 94633 -2093
rect 94911 -2371 94927 -2093
rect 94617 -2867 94927 -2371
rect 96477 349307 96787 355021
rect 105477 355779 105787 355795
rect 105477 355501 105493 355779
rect 105771 355501 105787 355779
rect 103617 354819 103927 354835
rect 103617 354541 103633 354819
rect 103911 354541 103927 354819
rect 101757 353859 102067 353875
rect 101757 353581 101773 353859
rect 102051 353581 102067 353859
rect 96477 349029 96493 349307
rect 96771 349029 96787 349307
rect 96477 331307 96787 349029
rect 96477 331029 96493 331307
rect 96771 331029 96787 331307
rect 96477 313307 96787 331029
rect 96477 313029 96493 313307
rect 96771 313029 96787 313307
rect 96477 295307 96787 313029
rect 96477 295029 96493 295307
rect 96771 295029 96787 295307
rect 96477 277307 96787 295029
rect 96477 277029 96493 277307
rect 96771 277029 96787 277307
rect 96477 259307 96787 277029
rect 96477 259029 96493 259307
rect 96771 259029 96787 259307
rect 96477 241307 96787 259029
rect 96477 241029 96493 241307
rect 96771 241029 96787 241307
rect 96477 223307 96787 241029
rect 96477 223029 96493 223307
rect 96771 223029 96787 223307
rect 96477 205307 96787 223029
rect 96477 205029 96493 205307
rect 96771 205029 96787 205307
rect 96477 187307 96787 205029
rect 96477 187029 96493 187307
rect 96771 187029 96787 187307
rect 96477 169307 96787 187029
rect 96477 169029 96493 169307
rect 96771 169029 96787 169307
rect 96477 151307 96787 169029
rect 96477 151029 96493 151307
rect 96771 151029 96787 151307
rect 96477 133307 96787 151029
rect 96477 133029 96493 133307
rect 96771 133029 96787 133307
rect 96477 115307 96787 133029
rect 96477 115029 96493 115307
rect 96771 115029 96787 115307
rect 96477 97307 96787 115029
rect 96477 97029 96493 97307
rect 96771 97029 96787 97307
rect 96477 79307 96787 97029
rect 96477 79029 96493 79307
rect 96771 79029 96787 79307
rect 96477 61307 96787 79029
rect 96477 61029 96493 61307
rect 96771 61029 96787 61307
rect 96477 43307 96787 61029
rect 96477 43029 96493 43307
rect 96771 43029 96787 43307
rect 96477 25307 96787 43029
rect 96477 25029 96493 25307
rect 96771 25029 96787 25307
rect 96477 7307 96787 25029
rect 96477 7029 96493 7307
rect 96771 7029 96787 7307
rect 87477 -3811 87493 -3533
rect 87771 -3811 87787 -3533
rect 87477 -3827 87787 -3811
rect 96477 -3053 96787 7029
rect 99897 352899 100207 352915
rect 99897 352621 99913 352899
rect 100191 352621 100207 352899
rect 99897 334727 100207 352621
rect 99897 334449 99913 334727
rect 100191 334449 100207 334727
rect 99897 316727 100207 334449
rect 99897 316449 99913 316727
rect 100191 316449 100207 316727
rect 99897 298727 100207 316449
rect 99897 298449 99913 298727
rect 100191 298449 100207 298727
rect 99897 280727 100207 298449
rect 99897 280449 99913 280727
rect 100191 280449 100207 280727
rect 99897 262727 100207 280449
rect 99897 262449 99913 262727
rect 100191 262449 100207 262727
rect 99897 244727 100207 262449
rect 99897 244449 99913 244727
rect 100191 244449 100207 244727
rect 99897 226727 100207 244449
rect 99897 226449 99913 226727
rect 100191 226449 100207 226727
rect 99897 208727 100207 226449
rect 99897 208449 99913 208727
rect 100191 208449 100207 208727
rect 99897 190727 100207 208449
rect 99897 190449 99913 190727
rect 100191 190449 100207 190727
rect 99897 172727 100207 190449
rect 99897 172449 99913 172727
rect 100191 172449 100207 172727
rect 99897 154727 100207 172449
rect 99897 154449 99913 154727
rect 100191 154449 100207 154727
rect 99897 136727 100207 154449
rect 99897 136449 99913 136727
rect 100191 136449 100207 136727
rect 99897 118727 100207 136449
rect 99897 118449 99913 118727
rect 100191 118449 100207 118727
rect 99897 100727 100207 118449
rect 99897 100449 99913 100727
rect 100191 100449 100207 100727
rect 99897 82727 100207 100449
rect 99897 82449 99913 82727
rect 100191 82449 100207 82727
rect 99897 64727 100207 82449
rect 99897 64449 99913 64727
rect 100191 64449 100207 64727
rect 99897 46727 100207 64449
rect 99897 46449 99913 46727
rect 100191 46449 100207 46727
rect 99897 28727 100207 46449
rect 99897 28449 99913 28727
rect 100191 28449 100207 28727
rect 99897 10727 100207 28449
rect 99897 10449 99913 10727
rect 100191 10449 100207 10727
rect 99897 -653 100207 10449
rect 99897 -931 99913 -653
rect 100191 -931 100207 -653
rect 99897 -947 100207 -931
rect 101757 336587 102067 353581
rect 101757 336309 101773 336587
rect 102051 336309 102067 336587
rect 101757 318587 102067 336309
rect 101757 318309 101773 318587
rect 102051 318309 102067 318587
rect 101757 300587 102067 318309
rect 101757 300309 101773 300587
rect 102051 300309 102067 300587
rect 101757 282587 102067 300309
rect 101757 282309 101773 282587
rect 102051 282309 102067 282587
rect 101757 264587 102067 282309
rect 101757 264309 101773 264587
rect 102051 264309 102067 264587
rect 101757 246587 102067 264309
rect 101757 246309 101773 246587
rect 102051 246309 102067 246587
rect 101757 228587 102067 246309
rect 101757 228309 101773 228587
rect 102051 228309 102067 228587
rect 101757 210587 102067 228309
rect 101757 210309 101773 210587
rect 102051 210309 102067 210587
rect 101757 192587 102067 210309
rect 101757 192309 101773 192587
rect 102051 192309 102067 192587
rect 101757 174587 102067 192309
rect 101757 174309 101773 174587
rect 102051 174309 102067 174587
rect 101757 156587 102067 174309
rect 101757 156309 101773 156587
rect 102051 156309 102067 156587
rect 101757 138587 102067 156309
rect 101757 138309 101773 138587
rect 102051 138309 102067 138587
rect 101757 120587 102067 138309
rect 101757 120309 101773 120587
rect 102051 120309 102067 120587
rect 101757 102587 102067 120309
rect 101757 102309 101773 102587
rect 102051 102309 102067 102587
rect 101757 84587 102067 102309
rect 101757 84309 101773 84587
rect 102051 84309 102067 84587
rect 101757 66587 102067 84309
rect 101757 66309 101773 66587
rect 102051 66309 102067 66587
rect 101757 48587 102067 66309
rect 101757 48309 101773 48587
rect 102051 48309 102067 48587
rect 101757 30587 102067 48309
rect 101757 30309 101773 30587
rect 102051 30309 102067 30587
rect 101757 12587 102067 30309
rect 101757 12309 101773 12587
rect 102051 12309 102067 12587
rect 101757 -1613 102067 12309
rect 101757 -1891 101773 -1613
rect 102051 -1891 102067 -1613
rect 101757 -1907 102067 -1891
rect 103617 338447 103927 354541
rect 103617 338169 103633 338447
rect 103911 338169 103927 338447
rect 103617 320447 103927 338169
rect 103617 320169 103633 320447
rect 103911 320169 103927 320447
rect 103617 302447 103927 320169
rect 103617 302169 103633 302447
rect 103911 302169 103927 302447
rect 103617 284447 103927 302169
rect 103617 284169 103633 284447
rect 103911 284169 103927 284447
rect 103617 266447 103927 284169
rect 103617 266169 103633 266447
rect 103911 266169 103927 266447
rect 103617 248447 103927 266169
rect 103617 248169 103633 248447
rect 103911 248169 103927 248447
rect 103617 230447 103927 248169
rect 103617 230169 103633 230447
rect 103911 230169 103927 230447
rect 103617 212447 103927 230169
rect 103617 212169 103633 212447
rect 103911 212169 103927 212447
rect 103617 194447 103927 212169
rect 103617 194169 103633 194447
rect 103911 194169 103927 194447
rect 103617 176447 103927 194169
rect 103617 176169 103633 176447
rect 103911 176169 103927 176447
rect 103617 158447 103927 176169
rect 103617 158169 103633 158447
rect 103911 158169 103927 158447
rect 103617 140447 103927 158169
rect 103617 140169 103633 140447
rect 103911 140169 103927 140447
rect 103617 122447 103927 140169
rect 103617 122169 103633 122447
rect 103911 122169 103927 122447
rect 103617 104447 103927 122169
rect 103617 104169 103633 104447
rect 103911 104169 103927 104447
rect 103617 86447 103927 104169
rect 103617 86169 103633 86447
rect 103911 86169 103927 86447
rect 103617 68447 103927 86169
rect 103617 68169 103633 68447
rect 103911 68169 103927 68447
rect 103617 50447 103927 68169
rect 103617 50169 103633 50447
rect 103911 50169 103927 50447
rect 103617 32447 103927 50169
rect 103617 32169 103633 32447
rect 103911 32169 103927 32447
rect 103617 14447 103927 32169
rect 103617 14169 103633 14447
rect 103911 14169 103927 14447
rect 103617 -2573 103927 14169
rect 103617 -2851 103633 -2573
rect 103911 -2851 103927 -2573
rect 103617 -2867 103927 -2851
rect 105477 340307 105787 355501
rect 114477 355299 114787 355795
rect 114477 355021 114493 355299
rect 114771 355021 114787 355299
rect 112617 354339 112927 354835
rect 112617 354061 112633 354339
rect 112911 354061 112927 354339
rect 110757 353379 111067 353875
rect 110757 353101 110773 353379
rect 111051 353101 111067 353379
rect 105477 340029 105493 340307
rect 105771 340029 105787 340307
rect 105477 322307 105787 340029
rect 105477 322029 105493 322307
rect 105771 322029 105787 322307
rect 105477 304307 105787 322029
rect 105477 304029 105493 304307
rect 105771 304029 105787 304307
rect 105477 286307 105787 304029
rect 105477 286029 105493 286307
rect 105771 286029 105787 286307
rect 105477 268307 105787 286029
rect 105477 268029 105493 268307
rect 105771 268029 105787 268307
rect 105477 250307 105787 268029
rect 105477 250029 105493 250307
rect 105771 250029 105787 250307
rect 105477 232307 105787 250029
rect 105477 232029 105493 232307
rect 105771 232029 105787 232307
rect 105477 214307 105787 232029
rect 105477 214029 105493 214307
rect 105771 214029 105787 214307
rect 105477 196307 105787 214029
rect 105477 196029 105493 196307
rect 105771 196029 105787 196307
rect 105477 178307 105787 196029
rect 105477 178029 105493 178307
rect 105771 178029 105787 178307
rect 105477 160307 105787 178029
rect 105477 160029 105493 160307
rect 105771 160029 105787 160307
rect 105477 142307 105787 160029
rect 105477 142029 105493 142307
rect 105771 142029 105787 142307
rect 105477 124307 105787 142029
rect 105477 124029 105493 124307
rect 105771 124029 105787 124307
rect 105477 106307 105787 124029
rect 105477 106029 105493 106307
rect 105771 106029 105787 106307
rect 105477 88307 105787 106029
rect 105477 88029 105493 88307
rect 105771 88029 105787 88307
rect 105477 70307 105787 88029
rect 105477 70029 105493 70307
rect 105771 70029 105787 70307
rect 105477 52307 105787 70029
rect 105477 52029 105493 52307
rect 105771 52029 105787 52307
rect 105477 34307 105787 52029
rect 105477 34029 105493 34307
rect 105771 34029 105787 34307
rect 105477 16307 105787 34029
rect 105477 16029 105493 16307
rect 105771 16029 105787 16307
rect 96477 -3331 96493 -3053
rect 96771 -3331 96787 -3053
rect 96477 -3827 96787 -3331
rect 105477 -3533 105787 16029
rect 108897 352419 109207 352915
rect 108897 352141 108913 352419
rect 109191 352141 109207 352419
rect 108897 343727 109207 352141
rect 108897 343449 108913 343727
rect 109191 343449 109207 343727
rect 108897 325727 109207 343449
rect 108897 325449 108913 325727
rect 109191 325449 109207 325727
rect 108897 307727 109207 325449
rect 108897 307449 108913 307727
rect 109191 307449 109207 307727
rect 108897 289727 109207 307449
rect 108897 289449 108913 289727
rect 109191 289449 109207 289727
rect 108897 271727 109207 289449
rect 108897 271449 108913 271727
rect 109191 271449 109207 271727
rect 108897 253727 109207 271449
rect 108897 253449 108913 253727
rect 109191 253449 109207 253727
rect 108897 235727 109207 253449
rect 108897 235449 108913 235727
rect 109191 235449 109207 235727
rect 108897 217727 109207 235449
rect 108897 217449 108913 217727
rect 109191 217449 109207 217727
rect 108897 199727 109207 217449
rect 108897 199449 108913 199727
rect 109191 199449 109207 199727
rect 108897 181727 109207 199449
rect 108897 181449 108913 181727
rect 109191 181449 109207 181727
rect 108897 163727 109207 181449
rect 108897 163449 108913 163727
rect 109191 163449 109207 163727
rect 108897 145727 109207 163449
rect 108897 145449 108913 145727
rect 109191 145449 109207 145727
rect 108897 127727 109207 145449
rect 108897 127449 108913 127727
rect 109191 127449 109207 127727
rect 108897 109727 109207 127449
rect 108897 109449 108913 109727
rect 109191 109449 109207 109727
rect 108897 91727 109207 109449
rect 108897 91449 108913 91727
rect 109191 91449 109207 91727
rect 108897 73727 109207 91449
rect 108897 73449 108913 73727
rect 109191 73449 109207 73727
rect 108897 55727 109207 73449
rect 108897 55449 108913 55727
rect 109191 55449 109207 55727
rect 108897 37727 109207 55449
rect 108897 37449 108913 37727
rect 109191 37449 109207 37727
rect 108897 19727 109207 37449
rect 108897 19449 108913 19727
rect 109191 19449 109207 19727
rect 108897 1727 109207 19449
rect 108897 1449 108913 1727
rect 109191 1449 109207 1727
rect 108897 -173 109207 1449
rect 108897 -451 108913 -173
rect 109191 -451 109207 -173
rect 108897 -947 109207 -451
rect 110757 345587 111067 353101
rect 110757 345309 110773 345587
rect 111051 345309 111067 345587
rect 110757 327587 111067 345309
rect 110757 327309 110773 327587
rect 111051 327309 111067 327587
rect 110757 309587 111067 327309
rect 110757 309309 110773 309587
rect 111051 309309 111067 309587
rect 110757 291587 111067 309309
rect 110757 291309 110773 291587
rect 111051 291309 111067 291587
rect 110757 273587 111067 291309
rect 110757 273309 110773 273587
rect 111051 273309 111067 273587
rect 110757 255587 111067 273309
rect 110757 255309 110773 255587
rect 111051 255309 111067 255587
rect 110757 237587 111067 255309
rect 110757 237309 110773 237587
rect 111051 237309 111067 237587
rect 110757 219587 111067 237309
rect 110757 219309 110773 219587
rect 111051 219309 111067 219587
rect 110757 201587 111067 219309
rect 110757 201309 110773 201587
rect 111051 201309 111067 201587
rect 110757 183587 111067 201309
rect 110757 183309 110773 183587
rect 111051 183309 111067 183587
rect 110757 165587 111067 183309
rect 110757 165309 110773 165587
rect 111051 165309 111067 165587
rect 110757 147587 111067 165309
rect 110757 147309 110773 147587
rect 111051 147309 111067 147587
rect 110757 129587 111067 147309
rect 110757 129309 110773 129587
rect 111051 129309 111067 129587
rect 110757 111587 111067 129309
rect 110757 111309 110773 111587
rect 111051 111309 111067 111587
rect 110757 93587 111067 111309
rect 110757 93309 110773 93587
rect 111051 93309 111067 93587
rect 110757 75587 111067 93309
rect 110757 75309 110773 75587
rect 111051 75309 111067 75587
rect 110757 57587 111067 75309
rect 110757 57309 110773 57587
rect 111051 57309 111067 57587
rect 110757 39587 111067 57309
rect 110757 39309 110773 39587
rect 111051 39309 111067 39587
rect 110757 21587 111067 39309
rect 110757 21309 110773 21587
rect 111051 21309 111067 21587
rect 110757 3587 111067 21309
rect 110757 3309 110773 3587
rect 111051 3309 111067 3587
rect 110757 -1133 111067 3309
rect 110757 -1411 110773 -1133
rect 111051 -1411 111067 -1133
rect 110757 -1907 111067 -1411
rect 112617 347447 112927 354061
rect 112617 347169 112633 347447
rect 112911 347169 112927 347447
rect 112617 329447 112927 347169
rect 112617 329169 112633 329447
rect 112911 329169 112927 329447
rect 112617 311447 112927 329169
rect 112617 311169 112633 311447
rect 112911 311169 112927 311447
rect 112617 293447 112927 311169
rect 112617 293169 112633 293447
rect 112911 293169 112927 293447
rect 112617 275447 112927 293169
rect 112617 275169 112633 275447
rect 112911 275169 112927 275447
rect 112617 257447 112927 275169
rect 112617 257169 112633 257447
rect 112911 257169 112927 257447
rect 112617 239447 112927 257169
rect 112617 239169 112633 239447
rect 112911 239169 112927 239447
rect 112617 221447 112927 239169
rect 112617 221169 112633 221447
rect 112911 221169 112927 221447
rect 112617 203447 112927 221169
rect 112617 203169 112633 203447
rect 112911 203169 112927 203447
rect 112617 185447 112927 203169
rect 112617 185169 112633 185447
rect 112911 185169 112927 185447
rect 112617 167447 112927 185169
rect 112617 167169 112633 167447
rect 112911 167169 112927 167447
rect 112617 149447 112927 167169
rect 112617 149169 112633 149447
rect 112911 149169 112927 149447
rect 112617 131447 112927 149169
rect 112617 131169 112633 131447
rect 112911 131169 112927 131447
rect 112617 113447 112927 131169
rect 112617 113169 112633 113447
rect 112911 113169 112927 113447
rect 112617 95447 112927 113169
rect 112617 95169 112633 95447
rect 112911 95169 112927 95447
rect 112617 77447 112927 95169
rect 112617 77169 112633 77447
rect 112911 77169 112927 77447
rect 112617 59447 112927 77169
rect 112617 59169 112633 59447
rect 112911 59169 112927 59447
rect 112617 41447 112927 59169
rect 112617 41169 112633 41447
rect 112911 41169 112927 41447
rect 112617 23447 112927 41169
rect 112617 23169 112633 23447
rect 112911 23169 112927 23447
rect 112617 5447 112927 23169
rect 112617 5169 112633 5447
rect 112911 5169 112927 5447
rect 112617 -2093 112927 5169
rect 112617 -2371 112633 -2093
rect 112911 -2371 112927 -2093
rect 112617 -2867 112927 -2371
rect 114477 349307 114787 355021
rect 123477 355779 123787 355795
rect 123477 355501 123493 355779
rect 123771 355501 123787 355779
rect 121617 354819 121927 354835
rect 121617 354541 121633 354819
rect 121911 354541 121927 354819
rect 119757 353859 120067 353875
rect 119757 353581 119773 353859
rect 120051 353581 120067 353859
rect 114477 349029 114493 349307
rect 114771 349029 114787 349307
rect 114477 331307 114787 349029
rect 114477 331029 114493 331307
rect 114771 331029 114787 331307
rect 114477 313307 114787 331029
rect 114477 313029 114493 313307
rect 114771 313029 114787 313307
rect 114477 295307 114787 313029
rect 114477 295029 114493 295307
rect 114771 295029 114787 295307
rect 114477 277307 114787 295029
rect 114477 277029 114493 277307
rect 114771 277029 114787 277307
rect 114477 259307 114787 277029
rect 114477 259029 114493 259307
rect 114771 259029 114787 259307
rect 114477 241307 114787 259029
rect 114477 241029 114493 241307
rect 114771 241029 114787 241307
rect 114477 223307 114787 241029
rect 114477 223029 114493 223307
rect 114771 223029 114787 223307
rect 114477 205307 114787 223029
rect 114477 205029 114493 205307
rect 114771 205029 114787 205307
rect 114477 187307 114787 205029
rect 114477 187029 114493 187307
rect 114771 187029 114787 187307
rect 114477 169307 114787 187029
rect 114477 169029 114493 169307
rect 114771 169029 114787 169307
rect 114477 151307 114787 169029
rect 114477 151029 114493 151307
rect 114771 151029 114787 151307
rect 114477 133307 114787 151029
rect 114477 133029 114493 133307
rect 114771 133029 114787 133307
rect 114477 115307 114787 133029
rect 114477 115029 114493 115307
rect 114771 115029 114787 115307
rect 114477 97307 114787 115029
rect 114477 97029 114493 97307
rect 114771 97029 114787 97307
rect 114477 79307 114787 97029
rect 114477 79029 114493 79307
rect 114771 79029 114787 79307
rect 114477 61307 114787 79029
rect 114477 61029 114493 61307
rect 114771 61029 114787 61307
rect 114477 43307 114787 61029
rect 114477 43029 114493 43307
rect 114771 43029 114787 43307
rect 114477 25307 114787 43029
rect 114477 25029 114493 25307
rect 114771 25029 114787 25307
rect 114477 7307 114787 25029
rect 114477 7029 114493 7307
rect 114771 7029 114787 7307
rect 105477 -3811 105493 -3533
rect 105771 -3811 105787 -3533
rect 105477 -3827 105787 -3811
rect 114477 -3053 114787 7029
rect 117897 352899 118207 352915
rect 117897 352621 117913 352899
rect 118191 352621 118207 352899
rect 117897 334727 118207 352621
rect 117897 334449 117913 334727
rect 118191 334449 118207 334727
rect 117897 316727 118207 334449
rect 117897 316449 117913 316727
rect 118191 316449 118207 316727
rect 117897 298727 118207 316449
rect 117897 298449 117913 298727
rect 118191 298449 118207 298727
rect 117897 280727 118207 298449
rect 117897 280449 117913 280727
rect 118191 280449 118207 280727
rect 117897 262727 118207 280449
rect 117897 262449 117913 262727
rect 118191 262449 118207 262727
rect 117897 244727 118207 262449
rect 117897 244449 117913 244727
rect 118191 244449 118207 244727
rect 117897 226727 118207 244449
rect 117897 226449 117913 226727
rect 118191 226449 118207 226727
rect 117897 208727 118207 226449
rect 117897 208449 117913 208727
rect 118191 208449 118207 208727
rect 117897 190727 118207 208449
rect 117897 190449 117913 190727
rect 118191 190449 118207 190727
rect 117897 172727 118207 190449
rect 117897 172449 117913 172727
rect 118191 172449 118207 172727
rect 117897 154727 118207 172449
rect 117897 154449 117913 154727
rect 118191 154449 118207 154727
rect 117897 136727 118207 154449
rect 117897 136449 117913 136727
rect 118191 136449 118207 136727
rect 117897 118727 118207 136449
rect 117897 118449 117913 118727
rect 118191 118449 118207 118727
rect 117897 100727 118207 118449
rect 117897 100449 117913 100727
rect 118191 100449 118207 100727
rect 117897 82727 118207 100449
rect 117897 82449 117913 82727
rect 118191 82449 118207 82727
rect 117897 64727 118207 82449
rect 117897 64449 117913 64727
rect 118191 64449 118207 64727
rect 117897 46727 118207 64449
rect 117897 46449 117913 46727
rect 118191 46449 118207 46727
rect 117897 28727 118207 46449
rect 117897 28449 117913 28727
rect 118191 28449 118207 28727
rect 117897 10727 118207 28449
rect 117897 10449 117913 10727
rect 118191 10449 118207 10727
rect 117897 -653 118207 10449
rect 117897 -931 117913 -653
rect 118191 -931 118207 -653
rect 117897 -947 118207 -931
rect 119757 336587 120067 353581
rect 119757 336309 119773 336587
rect 120051 336309 120067 336587
rect 119757 318587 120067 336309
rect 119757 318309 119773 318587
rect 120051 318309 120067 318587
rect 119757 300587 120067 318309
rect 119757 300309 119773 300587
rect 120051 300309 120067 300587
rect 119757 282587 120067 300309
rect 119757 282309 119773 282587
rect 120051 282309 120067 282587
rect 119757 264587 120067 282309
rect 119757 264309 119773 264587
rect 120051 264309 120067 264587
rect 119757 246587 120067 264309
rect 119757 246309 119773 246587
rect 120051 246309 120067 246587
rect 119757 228587 120067 246309
rect 119757 228309 119773 228587
rect 120051 228309 120067 228587
rect 119757 210587 120067 228309
rect 119757 210309 119773 210587
rect 120051 210309 120067 210587
rect 119757 192587 120067 210309
rect 119757 192309 119773 192587
rect 120051 192309 120067 192587
rect 119757 174587 120067 192309
rect 119757 174309 119773 174587
rect 120051 174309 120067 174587
rect 119757 156587 120067 174309
rect 119757 156309 119773 156587
rect 120051 156309 120067 156587
rect 119757 138587 120067 156309
rect 119757 138309 119773 138587
rect 120051 138309 120067 138587
rect 119757 120587 120067 138309
rect 119757 120309 119773 120587
rect 120051 120309 120067 120587
rect 119757 102587 120067 120309
rect 119757 102309 119773 102587
rect 120051 102309 120067 102587
rect 119757 84587 120067 102309
rect 119757 84309 119773 84587
rect 120051 84309 120067 84587
rect 119757 66587 120067 84309
rect 119757 66309 119773 66587
rect 120051 66309 120067 66587
rect 119757 48587 120067 66309
rect 119757 48309 119773 48587
rect 120051 48309 120067 48587
rect 119757 30587 120067 48309
rect 119757 30309 119773 30587
rect 120051 30309 120067 30587
rect 119757 12587 120067 30309
rect 119757 12309 119773 12587
rect 120051 12309 120067 12587
rect 119757 -1613 120067 12309
rect 119757 -1891 119773 -1613
rect 120051 -1891 120067 -1613
rect 119757 -1907 120067 -1891
rect 121617 338447 121927 354541
rect 121617 338169 121633 338447
rect 121911 338169 121927 338447
rect 121617 320447 121927 338169
rect 121617 320169 121633 320447
rect 121911 320169 121927 320447
rect 121617 302447 121927 320169
rect 121617 302169 121633 302447
rect 121911 302169 121927 302447
rect 121617 284447 121927 302169
rect 121617 284169 121633 284447
rect 121911 284169 121927 284447
rect 121617 266447 121927 284169
rect 121617 266169 121633 266447
rect 121911 266169 121927 266447
rect 121617 248447 121927 266169
rect 121617 248169 121633 248447
rect 121911 248169 121927 248447
rect 121617 230447 121927 248169
rect 121617 230169 121633 230447
rect 121911 230169 121927 230447
rect 121617 212447 121927 230169
rect 121617 212169 121633 212447
rect 121911 212169 121927 212447
rect 121617 194447 121927 212169
rect 121617 194169 121633 194447
rect 121911 194169 121927 194447
rect 121617 176447 121927 194169
rect 121617 176169 121633 176447
rect 121911 176169 121927 176447
rect 121617 158447 121927 176169
rect 121617 158169 121633 158447
rect 121911 158169 121927 158447
rect 121617 140447 121927 158169
rect 121617 140169 121633 140447
rect 121911 140169 121927 140447
rect 121617 122447 121927 140169
rect 121617 122169 121633 122447
rect 121911 122169 121927 122447
rect 121617 104447 121927 122169
rect 121617 104169 121633 104447
rect 121911 104169 121927 104447
rect 121617 86447 121927 104169
rect 121617 86169 121633 86447
rect 121911 86169 121927 86447
rect 121617 68447 121927 86169
rect 121617 68169 121633 68447
rect 121911 68169 121927 68447
rect 121617 50447 121927 68169
rect 121617 50169 121633 50447
rect 121911 50169 121927 50447
rect 121617 32447 121927 50169
rect 121617 32169 121633 32447
rect 121911 32169 121927 32447
rect 121617 14447 121927 32169
rect 121617 14169 121633 14447
rect 121911 14169 121927 14447
rect 121617 -2573 121927 14169
rect 121617 -2851 121633 -2573
rect 121911 -2851 121927 -2573
rect 121617 -2867 121927 -2851
rect 123477 340307 123787 355501
rect 132477 355299 132787 355795
rect 132477 355021 132493 355299
rect 132771 355021 132787 355299
rect 130617 354339 130927 354835
rect 130617 354061 130633 354339
rect 130911 354061 130927 354339
rect 128757 353379 129067 353875
rect 128757 353101 128773 353379
rect 129051 353101 129067 353379
rect 123477 340029 123493 340307
rect 123771 340029 123787 340307
rect 123477 322307 123787 340029
rect 123477 322029 123493 322307
rect 123771 322029 123787 322307
rect 123477 304307 123787 322029
rect 123477 304029 123493 304307
rect 123771 304029 123787 304307
rect 123477 286307 123787 304029
rect 123477 286029 123493 286307
rect 123771 286029 123787 286307
rect 123477 268307 123787 286029
rect 123477 268029 123493 268307
rect 123771 268029 123787 268307
rect 123477 250307 123787 268029
rect 123477 250029 123493 250307
rect 123771 250029 123787 250307
rect 123477 232307 123787 250029
rect 123477 232029 123493 232307
rect 123771 232029 123787 232307
rect 123477 214307 123787 232029
rect 123477 214029 123493 214307
rect 123771 214029 123787 214307
rect 123477 196307 123787 214029
rect 123477 196029 123493 196307
rect 123771 196029 123787 196307
rect 123477 178307 123787 196029
rect 123477 178029 123493 178307
rect 123771 178029 123787 178307
rect 123477 160307 123787 178029
rect 123477 160029 123493 160307
rect 123771 160029 123787 160307
rect 123477 142307 123787 160029
rect 123477 142029 123493 142307
rect 123771 142029 123787 142307
rect 123477 124307 123787 142029
rect 123477 124029 123493 124307
rect 123771 124029 123787 124307
rect 123477 106307 123787 124029
rect 123477 106029 123493 106307
rect 123771 106029 123787 106307
rect 123477 88307 123787 106029
rect 123477 88029 123493 88307
rect 123771 88029 123787 88307
rect 123477 70307 123787 88029
rect 123477 70029 123493 70307
rect 123771 70029 123787 70307
rect 123477 52307 123787 70029
rect 123477 52029 123493 52307
rect 123771 52029 123787 52307
rect 123477 34307 123787 52029
rect 123477 34029 123493 34307
rect 123771 34029 123787 34307
rect 123477 16307 123787 34029
rect 123477 16029 123493 16307
rect 123771 16029 123787 16307
rect 114477 -3331 114493 -3053
rect 114771 -3331 114787 -3053
rect 114477 -3827 114787 -3331
rect 123477 -3533 123787 16029
rect 126897 352419 127207 352915
rect 126897 352141 126913 352419
rect 127191 352141 127207 352419
rect 126897 343727 127207 352141
rect 126897 343449 126913 343727
rect 127191 343449 127207 343727
rect 126897 325727 127207 343449
rect 126897 325449 126913 325727
rect 127191 325449 127207 325727
rect 126897 307727 127207 325449
rect 126897 307449 126913 307727
rect 127191 307449 127207 307727
rect 126897 289727 127207 307449
rect 126897 289449 126913 289727
rect 127191 289449 127207 289727
rect 126897 271727 127207 289449
rect 126897 271449 126913 271727
rect 127191 271449 127207 271727
rect 126897 253727 127207 271449
rect 126897 253449 126913 253727
rect 127191 253449 127207 253727
rect 126897 235727 127207 253449
rect 126897 235449 126913 235727
rect 127191 235449 127207 235727
rect 126897 217727 127207 235449
rect 126897 217449 126913 217727
rect 127191 217449 127207 217727
rect 126897 199727 127207 217449
rect 126897 199449 126913 199727
rect 127191 199449 127207 199727
rect 126897 181727 127207 199449
rect 126897 181449 126913 181727
rect 127191 181449 127207 181727
rect 126897 163727 127207 181449
rect 126897 163449 126913 163727
rect 127191 163449 127207 163727
rect 126897 145727 127207 163449
rect 126897 145449 126913 145727
rect 127191 145449 127207 145727
rect 126897 127727 127207 145449
rect 126897 127449 126913 127727
rect 127191 127449 127207 127727
rect 126897 109727 127207 127449
rect 126897 109449 126913 109727
rect 127191 109449 127207 109727
rect 126897 91727 127207 109449
rect 126897 91449 126913 91727
rect 127191 91449 127207 91727
rect 126897 73727 127207 91449
rect 126897 73449 126913 73727
rect 127191 73449 127207 73727
rect 126897 55727 127207 73449
rect 126897 55449 126913 55727
rect 127191 55449 127207 55727
rect 126897 37727 127207 55449
rect 126897 37449 126913 37727
rect 127191 37449 127207 37727
rect 126897 19727 127207 37449
rect 126897 19449 126913 19727
rect 127191 19449 127207 19727
rect 126897 1727 127207 19449
rect 126897 1449 126913 1727
rect 127191 1449 127207 1727
rect 126897 -173 127207 1449
rect 126897 -451 126913 -173
rect 127191 -451 127207 -173
rect 126897 -947 127207 -451
rect 128757 345587 129067 353101
rect 128757 345309 128773 345587
rect 129051 345309 129067 345587
rect 128757 327587 129067 345309
rect 128757 327309 128773 327587
rect 129051 327309 129067 327587
rect 128757 309587 129067 327309
rect 128757 309309 128773 309587
rect 129051 309309 129067 309587
rect 128757 291587 129067 309309
rect 128757 291309 128773 291587
rect 129051 291309 129067 291587
rect 128757 273587 129067 291309
rect 128757 273309 128773 273587
rect 129051 273309 129067 273587
rect 128757 255587 129067 273309
rect 128757 255309 128773 255587
rect 129051 255309 129067 255587
rect 128757 237587 129067 255309
rect 128757 237309 128773 237587
rect 129051 237309 129067 237587
rect 128757 219587 129067 237309
rect 128757 219309 128773 219587
rect 129051 219309 129067 219587
rect 128757 201587 129067 219309
rect 128757 201309 128773 201587
rect 129051 201309 129067 201587
rect 128757 183587 129067 201309
rect 128757 183309 128773 183587
rect 129051 183309 129067 183587
rect 128757 165587 129067 183309
rect 128757 165309 128773 165587
rect 129051 165309 129067 165587
rect 128757 147587 129067 165309
rect 128757 147309 128773 147587
rect 129051 147309 129067 147587
rect 128757 129587 129067 147309
rect 128757 129309 128773 129587
rect 129051 129309 129067 129587
rect 128757 111587 129067 129309
rect 128757 111309 128773 111587
rect 129051 111309 129067 111587
rect 128757 93587 129067 111309
rect 128757 93309 128773 93587
rect 129051 93309 129067 93587
rect 128757 75587 129067 93309
rect 128757 75309 128773 75587
rect 129051 75309 129067 75587
rect 128757 57587 129067 75309
rect 128757 57309 128773 57587
rect 129051 57309 129067 57587
rect 128757 39587 129067 57309
rect 128757 39309 128773 39587
rect 129051 39309 129067 39587
rect 128757 21587 129067 39309
rect 128757 21309 128773 21587
rect 129051 21309 129067 21587
rect 128757 3587 129067 21309
rect 128757 3309 128773 3587
rect 129051 3309 129067 3587
rect 128757 -1133 129067 3309
rect 128757 -1411 128773 -1133
rect 129051 -1411 129067 -1133
rect 128757 -1907 129067 -1411
rect 130617 347447 130927 354061
rect 130617 347169 130633 347447
rect 130911 347169 130927 347447
rect 130617 329447 130927 347169
rect 130617 329169 130633 329447
rect 130911 329169 130927 329447
rect 130617 311447 130927 329169
rect 130617 311169 130633 311447
rect 130911 311169 130927 311447
rect 130617 293447 130927 311169
rect 130617 293169 130633 293447
rect 130911 293169 130927 293447
rect 130617 275447 130927 293169
rect 130617 275169 130633 275447
rect 130911 275169 130927 275447
rect 130617 257447 130927 275169
rect 130617 257169 130633 257447
rect 130911 257169 130927 257447
rect 130617 239447 130927 257169
rect 130617 239169 130633 239447
rect 130911 239169 130927 239447
rect 130617 221447 130927 239169
rect 130617 221169 130633 221447
rect 130911 221169 130927 221447
rect 130617 203447 130927 221169
rect 130617 203169 130633 203447
rect 130911 203169 130927 203447
rect 130617 185447 130927 203169
rect 130617 185169 130633 185447
rect 130911 185169 130927 185447
rect 130617 167447 130927 185169
rect 130617 167169 130633 167447
rect 130911 167169 130927 167447
rect 130617 149447 130927 167169
rect 130617 149169 130633 149447
rect 130911 149169 130927 149447
rect 130617 131447 130927 149169
rect 130617 131169 130633 131447
rect 130911 131169 130927 131447
rect 130617 113447 130927 131169
rect 130617 113169 130633 113447
rect 130911 113169 130927 113447
rect 130617 95447 130927 113169
rect 130617 95169 130633 95447
rect 130911 95169 130927 95447
rect 130617 77447 130927 95169
rect 130617 77169 130633 77447
rect 130911 77169 130927 77447
rect 130617 59447 130927 77169
rect 130617 59169 130633 59447
rect 130911 59169 130927 59447
rect 130617 41447 130927 59169
rect 130617 41169 130633 41447
rect 130911 41169 130927 41447
rect 130617 23447 130927 41169
rect 130617 23169 130633 23447
rect 130911 23169 130927 23447
rect 130617 5447 130927 23169
rect 130617 5169 130633 5447
rect 130911 5169 130927 5447
rect 130617 -2093 130927 5169
rect 130617 -2371 130633 -2093
rect 130911 -2371 130927 -2093
rect 130617 -2867 130927 -2371
rect 132477 349307 132787 355021
rect 141477 355779 141787 355795
rect 141477 355501 141493 355779
rect 141771 355501 141787 355779
rect 139617 354819 139927 354835
rect 139617 354541 139633 354819
rect 139911 354541 139927 354819
rect 137757 353859 138067 353875
rect 137757 353581 137773 353859
rect 138051 353581 138067 353859
rect 132477 349029 132493 349307
rect 132771 349029 132787 349307
rect 132477 331307 132787 349029
rect 132477 331029 132493 331307
rect 132771 331029 132787 331307
rect 132477 313307 132787 331029
rect 132477 313029 132493 313307
rect 132771 313029 132787 313307
rect 132477 295307 132787 313029
rect 132477 295029 132493 295307
rect 132771 295029 132787 295307
rect 132477 277307 132787 295029
rect 132477 277029 132493 277307
rect 132771 277029 132787 277307
rect 132477 259307 132787 277029
rect 132477 259029 132493 259307
rect 132771 259029 132787 259307
rect 132477 241307 132787 259029
rect 132477 241029 132493 241307
rect 132771 241029 132787 241307
rect 132477 223307 132787 241029
rect 132477 223029 132493 223307
rect 132771 223029 132787 223307
rect 132477 205307 132787 223029
rect 132477 205029 132493 205307
rect 132771 205029 132787 205307
rect 132477 187307 132787 205029
rect 132477 187029 132493 187307
rect 132771 187029 132787 187307
rect 132477 169307 132787 187029
rect 132477 169029 132493 169307
rect 132771 169029 132787 169307
rect 132477 151307 132787 169029
rect 132477 151029 132493 151307
rect 132771 151029 132787 151307
rect 132477 133307 132787 151029
rect 132477 133029 132493 133307
rect 132771 133029 132787 133307
rect 132477 115307 132787 133029
rect 132477 115029 132493 115307
rect 132771 115029 132787 115307
rect 132477 97307 132787 115029
rect 132477 97029 132493 97307
rect 132771 97029 132787 97307
rect 132477 79307 132787 97029
rect 132477 79029 132493 79307
rect 132771 79029 132787 79307
rect 132477 61307 132787 79029
rect 132477 61029 132493 61307
rect 132771 61029 132787 61307
rect 132477 43307 132787 61029
rect 132477 43029 132493 43307
rect 132771 43029 132787 43307
rect 132477 25307 132787 43029
rect 132477 25029 132493 25307
rect 132771 25029 132787 25307
rect 132477 7307 132787 25029
rect 132477 7029 132493 7307
rect 132771 7029 132787 7307
rect 123477 -3811 123493 -3533
rect 123771 -3811 123787 -3533
rect 123477 -3827 123787 -3811
rect 132477 -3053 132787 7029
rect 135897 352899 136207 352915
rect 135897 352621 135913 352899
rect 136191 352621 136207 352899
rect 135897 334727 136207 352621
rect 135897 334449 135913 334727
rect 136191 334449 136207 334727
rect 135897 316727 136207 334449
rect 135897 316449 135913 316727
rect 136191 316449 136207 316727
rect 135897 298727 136207 316449
rect 135897 298449 135913 298727
rect 136191 298449 136207 298727
rect 135897 280727 136207 298449
rect 135897 280449 135913 280727
rect 136191 280449 136207 280727
rect 135897 262727 136207 280449
rect 135897 262449 135913 262727
rect 136191 262449 136207 262727
rect 135897 244727 136207 262449
rect 135897 244449 135913 244727
rect 136191 244449 136207 244727
rect 135897 226727 136207 244449
rect 135897 226449 135913 226727
rect 136191 226449 136207 226727
rect 135897 208727 136207 226449
rect 135897 208449 135913 208727
rect 136191 208449 136207 208727
rect 135897 190727 136207 208449
rect 135897 190449 135913 190727
rect 136191 190449 136207 190727
rect 135897 172727 136207 190449
rect 135897 172449 135913 172727
rect 136191 172449 136207 172727
rect 135897 154727 136207 172449
rect 135897 154449 135913 154727
rect 136191 154449 136207 154727
rect 135897 136727 136207 154449
rect 135897 136449 135913 136727
rect 136191 136449 136207 136727
rect 135897 118727 136207 136449
rect 135897 118449 135913 118727
rect 136191 118449 136207 118727
rect 135897 100727 136207 118449
rect 135897 100449 135913 100727
rect 136191 100449 136207 100727
rect 135897 82727 136207 100449
rect 135897 82449 135913 82727
rect 136191 82449 136207 82727
rect 135897 64727 136207 82449
rect 135897 64449 135913 64727
rect 136191 64449 136207 64727
rect 135897 46727 136207 64449
rect 135897 46449 135913 46727
rect 136191 46449 136207 46727
rect 135897 28727 136207 46449
rect 135897 28449 135913 28727
rect 136191 28449 136207 28727
rect 135897 10727 136207 28449
rect 135897 10449 135913 10727
rect 136191 10449 136207 10727
rect 135897 -653 136207 10449
rect 135897 -931 135913 -653
rect 136191 -931 136207 -653
rect 135897 -947 136207 -931
rect 137757 336587 138067 353581
rect 137757 336309 137773 336587
rect 138051 336309 138067 336587
rect 137757 318587 138067 336309
rect 137757 318309 137773 318587
rect 138051 318309 138067 318587
rect 137757 300587 138067 318309
rect 137757 300309 137773 300587
rect 138051 300309 138067 300587
rect 137757 282587 138067 300309
rect 137757 282309 137773 282587
rect 138051 282309 138067 282587
rect 137757 264587 138067 282309
rect 137757 264309 137773 264587
rect 138051 264309 138067 264587
rect 137757 246587 138067 264309
rect 137757 246309 137773 246587
rect 138051 246309 138067 246587
rect 137757 228587 138067 246309
rect 137757 228309 137773 228587
rect 138051 228309 138067 228587
rect 137757 210587 138067 228309
rect 137757 210309 137773 210587
rect 138051 210309 138067 210587
rect 137757 192587 138067 210309
rect 137757 192309 137773 192587
rect 138051 192309 138067 192587
rect 137757 174587 138067 192309
rect 137757 174309 137773 174587
rect 138051 174309 138067 174587
rect 137757 156587 138067 174309
rect 137757 156309 137773 156587
rect 138051 156309 138067 156587
rect 137757 138587 138067 156309
rect 137757 138309 137773 138587
rect 138051 138309 138067 138587
rect 137757 120587 138067 138309
rect 137757 120309 137773 120587
rect 138051 120309 138067 120587
rect 137757 102587 138067 120309
rect 137757 102309 137773 102587
rect 138051 102309 138067 102587
rect 137757 84587 138067 102309
rect 137757 84309 137773 84587
rect 138051 84309 138067 84587
rect 137757 66587 138067 84309
rect 137757 66309 137773 66587
rect 138051 66309 138067 66587
rect 137757 48587 138067 66309
rect 137757 48309 137773 48587
rect 138051 48309 138067 48587
rect 137757 30587 138067 48309
rect 137757 30309 137773 30587
rect 138051 30309 138067 30587
rect 137757 12587 138067 30309
rect 137757 12309 137773 12587
rect 138051 12309 138067 12587
rect 137757 -1613 138067 12309
rect 137757 -1891 137773 -1613
rect 138051 -1891 138067 -1613
rect 137757 -1907 138067 -1891
rect 139617 338447 139927 354541
rect 139617 338169 139633 338447
rect 139911 338169 139927 338447
rect 139617 320447 139927 338169
rect 139617 320169 139633 320447
rect 139911 320169 139927 320447
rect 139617 302447 139927 320169
rect 139617 302169 139633 302447
rect 139911 302169 139927 302447
rect 139617 284447 139927 302169
rect 139617 284169 139633 284447
rect 139911 284169 139927 284447
rect 139617 266447 139927 284169
rect 139617 266169 139633 266447
rect 139911 266169 139927 266447
rect 139617 248447 139927 266169
rect 139617 248169 139633 248447
rect 139911 248169 139927 248447
rect 139617 230447 139927 248169
rect 139617 230169 139633 230447
rect 139911 230169 139927 230447
rect 139617 212447 139927 230169
rect 139617 212169 139633 212447
rect 139911 212169 139927 212447
rect 139617 194447 139927 212169
rect 139617 194169 139633 194447
rect 139911 194169 139927 194447
rect 139617 176447 139927 194169
rect 139617 176169 139633 176447
rect 139911 176169 139927 176447
rect 139617 158447 139927 176169
rect 139617 158169 139633 158447
rect 139911 158169 139927 158447
rect 139617 140447 139927 158169
rect 139617 140169 139633 140447
rect 139911 140169 139927 140447
rect 139617 122447 139927 140169
rect 139617 122169 139633 122447
rect 139911 122169 139927 122447
rect 139617 104447 139927 122169
rect 139617 104169 139633 104447
rect 139911 104169 139927 104447
rect 139617 86447 139927 104169
rect 139617 86169 139633 86447
rect 139911 86169 139927 86447
rect 139617 68447 139927 86169
rect 139617 68169 139633 68447
rect 139911 68169 139927 68447
rect 139617 50447 139927 68169
rect 139617 50169 139633 50447
rect 139911 50169 139927 50447
rect 139617 32447 139927 50169
rect 139617 32169 139633 32447
rect 139911 32169 139927 32447
rect 139617 14447 139927 32169
rect 139617 14169 139633 14447
rect 139911 14169 139927 14447
rect 139617 -2573 139927 14169
rect 139617 -2851 139633 -2573
rect 139911 -2851 139927 -2573
rect 139617 -2867 139927 -2851
rect 141477 340307 141787 355501
rect 150477 355299 150787 355795
rect 150477 355021 150493 355299
rect 150771 355021 150787 355299
rect 148617 354339 148927 354835
rect 148617 354061 148633 354339
rect 148911 354061 148927 354339
rect 146757 353379 147067 353875
rect 146757 353101 146773 353379
rect 147051 353101 147067 353379
rect 141477 340029 141493 340307
rect 141771 340029 141787 340307
rect 141477 322307 141787 340029
rect 141477 322029 141493 322307
rect 141771 322029 141787 322307
rect 141477 304307 141787 322029
rect 141477 304029 141493 304307
rect 141771 304029 141787 304307
rect 141477 286307 141787 304029
rect 141477 286029 141493 286307
rect 141771 286029 141787 286307
rect 141477 268307 141787 286029
rect 141477 268029 141493 268307
rect 141771 268029 141787 268307
rect 141477 250307 141787 268029
rect 141477 250029 141493 250307
rect 141771 250029 141787 250307
rect 141477 232307 141787 250029
rect 141477 232029 141493 232307
rect 141771 232029 141787 232307
rect 141477 214307 141787 232029
rect 141477 214029 141493 214307
rect 141771 214029 141787 214307
rect 141477 196307 141787 214029
rect 141477 196029 141493 196307
rect 141771 196029 141787 196307
rect 141477 178307 141787 196029
rect 141477 178029 141493 178307
rect 141771 178029 141787 178307
rect 141477 160307 141787 178029
rect 141477 160029 141493 160307
rect 141771 160029 141787 160307
rect 141477 142307 141787 160029
rect 141477 142029 141493 142307
rect 141771 142029 141787 142307
rect 141477 124307 141787 142029
rect 141477 124029 141493 124307
rect 141771 124029 141787 124307
rect 141477 106307 141787 124029
rect 141477 106029 141493 106307
rect 141771 106029 141787 106307
rect 141477 88307 141787 106029
rect 141477 88029 141493 88307
rect 141771 88029 141787 88307
rect 141477 70307 141787 88029
rect 141477 70029 141493 70307
rect 141771 70029 141787 70307
rect 141477 52307 141787 70029
rect 141477 52029 141493 52307
rect 141771 52029 141787 52307
rect 141477 34307 141787 52029
rect 141477 34029 141493 34307
rect 141771 34029 141787 34307
rect 141477 16307 141787 34029
rect 141477 16029 141493 16307
rect 141771 16029 141787 16307
rect 132477 -3331 132493 -3053
rect 132771 -3331 132787 -3053
rect 132477 -3827 132787 -3331
rect 141477 -3533 141787 16029
rect 144897 352419 145207 352915
rect 144897 352141 144913 352419
rect 145191 352141 145207 352419
rect 144897 343727 145207 352141
rect 144897 343449 144913 343727
rect 145191 343449 145207 343727
rect 144897 325727 145207 343449
rect 144897 325449 144913 325727
rect 145191 325449 145207 325727
rect 144897 307727 145207 325449
rect 144897 307449 144913 307727
rect 145191 307449 145207 307727
rect 144897 289727 145207 307449
rect 144897 289449 144913 289727
rect 145191 289449 145207 289727
rect 144897 271727 145207 289449
rect 144897 271449 144913 271727
rect 145191 271449 145207 271727
rect 144897 253727 145207 271449
rect 144897 253449 144913 253727
rect 145191 253449 145207 253727
rect 144897 235727 145207 253449
rect 144897 235449 144913 235727
rect 145191 235449 145207 235727
rect 144897 217727 145207 235449
rect 144897 217449 144913 217727
rect 145191 217449 145207 217727
rect 144897 199727 145207 217449
rect 144897 199449 144913 199727
rect 145191 199449 145207 199727
rect 144897 181727 145207 199449
rect 144897 181449 144913 181727
rect 145191 181449 145207 181727
rect 144897 163727 145207 181449
rect 144897 163449 144913 163727
rect 145191 163449 145207 163727
rect 144897 145727 145207 163449
rect 144897 145449 144913 145727
rect 145191 145449 145207 145727
rect 144897 127727 145207 145449
rect 144897 127449 144913 127727
rect 145191 127449 145207 127727
rect 144897 109727 145207 127449
rect 144897 109449 144913 109727
rect 145191 109449 145207 109727
rect 144897 91727 145207 109449
rect 144897 91449 144913 91727
rect 145191 91449 145207 91727
rect 144897 73727 145207 91449
rect 144897 73449 144913 73727
rect 145191 73449 145207 73727
rect 144897 55727 145207 73449
rect 144897 55449 144913 55727
rect 145191 55449 145207 55727
rect 144897 37727 145207 55449
rect 144897 37449 144913 37727
rect 145191 37449 145207 37727
rect 144897 19727 145207 37449
rect 144897 19449 144913 19727
rect 145191 19449 145207 19727
rect 144897 1727 145207 19449
rect 144897 1449 144913 1727
rect 145191 1449 145207 1727
rect 144897 -173 145207 1449
rect 144897 -451 144913 -173
rect 145191 -451 145207 -173
rect 144897 -947 145207 -451
rect 146757 345587 147067 353101
rect 146757 345309 146773 345587
rect 147051 345309 147067 345587
rect 146757 327587 147067 345309
rect 146757 327309 146773 327587
rect 147051 327309 147067 327587
rect 146757 309587 147067 327309
rect 146757 309309 146773 309587
rect 147051 309309 147067 309587
rect 146757 291587 147067 309309
rect 146757 291309 146773 291587
rect 147051 291309 147067 291587
rect 146757 273587 147067 291309
rect 146757 273309 146773 273587
rect 147051 273309 147067 273587
rect 146757 255587 147067 273309
rect 146757 255309 146773 255587
rect 147051 255309 147067 255587
rect 146757 237587 147067 255309
rect 146757 237309 146773 237587
rect 147051 237309 147067 237587
rect 146757 219587 147067 237309
rect 146757 219309 146773 219587
rect 147051 219309 147067 219587
rect 146757 201587 147067 219309
rect 146757 201309 146773 201587
rect 147051 201309 147067 201587
rect 146757 183587 147067 201309
rect 146757 183309 146773 183587
rect 147051 183309 147067 183587
rect 146757 165587 147067 183309
rect 146757 165309 146773 165587
rect 147051 165309 147067 165587
rect 146757 147587 147067 165309
rect 146757 147309 146773 147587
rect 147051 147309 147067 147587
rect 146757 129587 147067 147309
rect 146757 129309 146773 129587
rect 147051 129309 147067 129587
rect 146757 111587 147067 129309
rect 146757 111309 146773 111587
rect 147051 111309 147067 111587
rect 146757 93587 147067 111309
rect 146757 93309 146773 93587
rect 147051 93309 147067 93587
rect 146757 75587 147067 93309
rect 146757 75309 146773 75587
rect 147051 75309 147067 75587
rect 146757 57587 147067 75309
rect 146757 57309 146773 57587
rect 147051 57309 147067 57587
rect 146757 39587 147067 57309
rect 146757 39309 146773 39587
rect 147051 39309 147067 39587
rect 146757 21587 147067 39309
rect 146757 21309 146773 21587
rect 147051 21309 147067 21587
rect 146757 3587 147067 21309
rect 146757 3309 146773 3587
rect 147051 3309 147067 3587
rect 146757 -1133 147067 3309
rect 146757 -1411 146773 -1133
rect 147051 -1411 147067 -1133
rect 146757 -1907 147067 -1411
rect 148617 347447 148927 354061
rect 148617 347169 148633 347447
rect 148911 347169 148927 347447
rect 148617 329447 148927 347169
rect 148617 329169 148633 329447
rect 148911 329169 148927 329447
rect 148617 311447 148927 329169
rect 148617 311169 148633 311447
rect 148911 311169 148927 311447
rect 148617 293447 148927 311169
rect 148617 293169 148633 293447
rect 148911 293169 148927 293447
rect 148617 275447 148927 293169
rect 148617 275169 148633 275447
rect 148911 275169 148927 275447
rect 148617 257447 148927 275169
rect 148617 257169 148633 257447
rect 148911 257169 148927 257447
rect 148617 239447 148927 257169
rect 148617 239169 148633 239447
rect 148911 239169 148927 239447
rect 148617 221447 148927 239169
rect 148617 221169 148633 221447
rect 148911 221169 148927 221447
rect 148617 203447 148927 221169
rect 148617 203169 148633 203447
rect 148911 203169 148927 203447
rect 148617 185447 148927 203169
rect 148617 185169 148633 185447
rect 148911 185169 148927 185447
rect 148617 167447 148927 185169
rect 148617 167169 148633 167447
rect 148911 167169 148927 167447
rect 148617 149447 148927 167169
rect 148617 149169 148633 149447
rect 148911 149169 148927 149447
rect 148617 131447 148927 149169
rect 148617 131169 148633 131447
rect 148911 131169 148927 131447
rect 148617 113447 148927 131169
rect 148617 113169 148633 113447
rect 148911 113169 148927 113447
rect 148617 95447 148927 113169
rect 148617 95169 148633 95447
rect 148911 95169 148927 95447
rect 148617 77447 148927 95169
rect 148617 77169 148633 77447
rect 148911 77169 148927 77447
rect 148617 59447 148927 77169
rect 148617 59169 148633 59447
rect 148911 59169 148927 59447
rect 148617 41447 148927 59169
rect 148617 41169 148633 41447
rect 148911 41169 148927 41447
rect 148617 23447 148927 41169
rect 148617 23169 148633 23447
rect 148911 23169 148927 23447
rect 148617 5447 148927 23169
rect 148617 5169 148633 5447
rect 148911 5169 148927 5447
rect 148617 -2093 148927 5169
rect 148617 -2371 148633 -2093
rect 148911 -2371 148927 -2093
rect 148617 -2867 148927 -2371
rect 150477 349307 150787 355021
rect 159477 355779 159787 355795
rect 159477 355501 159493 355779
rect 159771 355501 159787 355779
rect 157617 354819 157927 354835
rect 157617 354541 157633 354819
rect 157911 354541 157927 354819
rect 155757 353859 156067 353875
rect 155757 353581 155773 353859
rect 156051 353581 156067 353859
rect 150477 349029 150493 349307
rect 150771 349029 150787 349307
rect 150477 331307 150787 349029
rect 150477 331029 150493 331307
rect 150771 331029 150787 331307
rect 150477 313307 150787 331029
rect 150477 313029 150493 313307
rect 150771 313029 150787 313307
rect 150477 295307 150787 313029
rect 150477 295029 150493 295307
rect 150771 295029 150787 295307
rect 150477 277307 150787 295029
rect 150477 277029 150493 277307
rect 150771 277029 150787 277307
rect 150477 259307 150787 277029
rect 150477 259029 150493 259307
rect 150771 259029 150787 259307
rect 150477 241307 150787 259029
rect 150477 241029 150493 241307
rect 150771 241029 150787 241307
rect 150477 223307 150787 241029
rect 150477 223029 150493 223307
rect 150771 223029 150787 223307
rect 150477 205307 150787 223029
rect 150477 205029 150493 205307
rect 150771 205029 150787 205307
rect 150477 187307 150787 205029
rect 150477 187029 150493 187307
rect 150771 187029 150787 187307
rect 150477 169307 150787 187029
rect 150477 169029 150493 169307
rect 150771 169029 150787 169307
rect 150477 151307 150787 169029
rect 150477 151029 150493 151307
rect 150771 151029 150787 151307
rect 150477 133307 150787 151029
rect 150477 133029 150493 133307
rect 150771 133029 150787 133307
rect 150477 115307 150787 133029
rect 150477 115029 150493 115307
rect 150771 115029 150787 115307
rect 150477 97307 150787 115029
rect 150477 97029 150493 97307
rect 150771 97029 150787 97307
rect 150477 79307 150787 97029
rect 150477 79029 150493 79307
rect 150771 79029 150787 79307
rect 150477 61307 150787 79029
rect 150477 61029 150493 61307
rect 150771 61029 150787 61307
rect 150477 43307 150787 61029
rect 150477 43029 150493 43307
rect 150771 43029 150787 43307
rect 150477 25307 150787 43029
rect 150477 25029 150493 25307
rect 150771 25029 150787 25307
rect 150477 7307 150787 25029
rect 150477 7029 150493 7307
rect 150771 7029 150787 7307
rect 141477 -3811 141493 -3533
rect 141771 -3811 141787 -3533
rect 141477 -3827 141787 -3811
rect 150477 -3053 150787 7029
rect 153897 352899 154207 352915
rect 153897 352621 153913 352899
rect 154191 352621 154207 352899
rect 153897 334727 154207 352621
rect 153897 334449 153913 334727
rect 154191 334449 154207 334727
rect 153897 316727 154207 334449
rect 153897 316449 153913 316727
rect 154191 316449 154207 316727
rect 153897 298727 154207 316449
rect 153897 298449 153913 298727
rect 154191 298449 154207 298727
rect 153897 280727 154207 298449
rect 153897 280449 153913 280727
rect 154191 280449 154207 280727
rect 153897 262727 154207 280449
rect 153897 262449 153913 262727
rect 154191 262449 154207 262727
rect 153897 244727 154207 262449
rect 153897 244449 153913 244727
rect 154191 244449 154207 244727
rect 153897 226727 154207 244449
rect 153897 226449 153913 226727
rect 154191 226449 154207 226727
rect 153897 208727 154207 226449
rect 153897 208449 153913 208727
rect 154191 208449 154207 208727
rect 153897 190727 154207 208449
rect 153897 190449 153913 190727
rect 154191 190449 154207 190727
rect 153897 172727 154207 190449
rect 153897 172449 153913 172727
rect 154191 172449 154207 172727
rect 153897 154727 154207 172449
rect 153897 154449 153913 154727
rect 154191 154449 154207 154727
rect 153897 136727 154207 154449
rect 153897 136449 153913 136727
rect 154191 136449 154207 136727
rect 153897 118727 154207 136449
rect 153897 118449 153913 118727
rect 154191 118449 154207 118727
rect 153897 100727 154207 118449
rect 153897 100449 153913 100727
rect 154191 100449 154207 100727
rect 153897 82727 154207 100449
rect 153897 82449 153913 82727
rect 154191 82449 154207 82727
rect 153897 64727 154207 82449
rect 153897 64449 153913 64727
rect 154191 64449 154207 64727
rect 153897 46727 154207 64449
rect 153897 46449 153913 46727
rect 154191 46449 154207 46727
rect 153897 28727 154207 46449
rect 153897 28449 153913 28727
rect 154191 28449 154207 28727
rect 153897 10727 154207 28449
rect 153897 10449 153913 10727
rect 154191 10449 154207 10727
rect 153897 -653 154207 10449
rect 153897 -931 153913 -653
rect 154191 -931 154207 -653
rect 153897 -947 154207 -931
rect 155757 336587 156067 353581
rect 155757 336309 155773 336587
rect 156051 336309 156067 336587
rect 155757 318587 156067 336309
rect 155757 318309 155773 318587
rect 156051 318309 156067 318587
rect 155757 300587 156067 318309
rect 155757 300309 155773 300587
rect 156051 300309 156067 300587
rect 155757 282587 156067 300309
rect 155757 282309 155773 282587
rect 156051 282309 156067 282587
rect 155757 264587 156067 282309
rect 155757 264309 155773 264587
rect 156051 264309 156067 264587
rect 155757 246587 156067 264309
rect 155757 246309 155773 246587
rect 156051 246309 156067 246587
rect 155757 228587 156067 246309
rect 155757 228309 155773 228587
rect 156051 228309 156067 228587
rect 155757 210587 156067 228309
rect 155757 210309 155773 210587
rect 156051 210309 156067 210587
rect 155757 192587 156067 210309
rect 155757 192309 155773 192587
rect 156051 192309 156067 192587
rect 155757 174587 156067 192309
rect 155757 174309 155773 174587
rect 156051 174309 156067 174587
rect 155757 156587 156067 174309
rect 155757 156309 155773 156587
rect 156051 156309 156067 156587
rect 155757 138587 156067 156309
rect 155757 138309 155773 138587
rect 156051 138309 156067 138587
rect 155757 120587 156067 138309
rect 155757 120309 155773 120587
rect 156051 120309 156067 120587
rect 155757 102587 156067 120309
rect 155757 102309 155773 102587
rect 156051 102309 156067 102587
rect 155757 84587 156067 102309
rect 155757 84309 155773 84587
rect 156051 84309 156067 84587
rect 155757 66587 156067 84309
rect 155757 66309 155773 66587
rect 156051 66309 156067 66587
rect 155757 48587 156067 66309
rect 155757 48309 155773 48587
rect 156051 48309 156067 48587
rect 155757 30587 156067 48309
rect 155757 30309 155773 30587
rect 156051 30309 156067 30587
rect 155757 12587 156067 30309
rect 155757 12309 155773 12587
rect 156051 12309 156067 12587
rect 155757 -1613 156067 12309
rect 155757 -1891 155773 -1613
rect 156051 -1891 156067 -1613
rect 155757 -1907 156067 -1891
rect 157617 338447 157927 354541
rect 157617 338169 157633 338447
rect 157911 338169 157927 338447
rect 157617 320447 157927 338169
rect 157617 320169 157633 320447
rect 157911 320169 157927 320447
rect 157617 302447 157927 320169
rect 157617 302169 157633 302447
rect 157911 302169 157927 302447
rect 157617 284447 157927 302169
rect 157617 284169 157633 284447
rect 157911 284169 157927 284447
rect 157617 266447 157927 284169
rect 157617 266169 157633 266447
rect 157911 266169 157927 266447
rect 157617 248447 157927 266169
rect 157617 248169 157633 248447
rect 157911 248169 157927 248447
rect 157617 230447 157927 248169
rect 157617 230169 157633 230447
rect 157911 230169 157927 230447
rect 157617 212447 157927 230169
rect 157617 212169 157633 212447
rect 157911 212169 157927 212447
rect 157617 194447 157927 212169
rect 157617 194169 157633 194447
rect 157911 194169 157927 194447
rect 157617 176447 157927 194169
rect 157617 176169 157633 176447
rect 157911 176169 157927 176447
rect 157617 158447 157927 176169
rect 157617 158169 157633 158447
rect 157911 158169 157927 158447
rect 157617 140447 157927 158169
rect 157617 140169 157633 140447
rect 157911 140169 157927 140447
rect 157617 122447 157927 140169
rect 157617 122169 157633 122447
rect 157911 122169 157927 122447
rect 157617 104447 157927 122169
rect 157617 104169 157633 104447
rect 157911 104169 157927 104447
rect 157617 86447 157927 104169
rect 157617 86169 157633 86447
rect 157911 86169 157927 86447
rect 157617 68447 157927 86169
rect 157617 68169 157633 68447
rect 157911 68169 157927 68447
rect 157617 50447 157927 68169
rect 157617 50169 157633 50447
rect 157911 50169 157927 50447
rect 157617 32447 157927 50169
rect 157617 32169 157633 32447
rect 157911 32169 157927 32447
rect 157617 14447 157927 32169
rect 157617 14169 157633 14447
rect 157911 14169 157927 14447
rect 157617 -2573 157927 14169
rect 157617 -2851 157633 -2573
rect 157911 -2851 157927 -2573
rect 157617 -2867 157927 -2851
rect 159477 340307 159787 355501
rect 168477 355299 168787 355795
rect 168477 355021 168493 355299
rect 168771 355021 168787 355299
rect 166617 354339 166927 354835
rect 166617 354061 166633 354339
rect 166911 354061 166927 354339
rect 164757 353379 165067 353875
rect 164757 353101 164773 353379
rect 165051 353101 165067 353379
rect 159477 340029 159493 340307
rect 159771 340029 159787 340307
rect 159477 322307 159787 340029
rect 159477 322029 159493 322307
rect 159771 322029 159787 322307
rect 159477 304307 159787 322029
rect 159477 304029 159493 304307
rect 159771 304029 159787 304307
rect 159477 286307 159787 304029
rect 159477 286029 159493 286307
rect 159771 286029 159787 286307
rect 159477 268307 159787 286029
rect 159477 268029 159493 268307
rect 159771 268029 159787 268307
rect 159477 250307 159787 268029
rect 159477 250029 159493 250307
rect 159771 250029 159787 250307
rect 159477 232307 159787 250029
rect 159477 232029 159493 232307
rect 159771 232029 159787 232307
rect 159477 214307 159787 232029
rect 159477 214029 159493 214307
rect 159771 214029 159787 214307
rect 159477 196307 159787 214029
rect 159477 196029 159493 196307
rect 159771 196029 159787 196307
rect 159477 178307 159787 196029
rect 159477 178029 159493 178307
rect 159771 178029 159787 178307
rect 159477 160307 159787 178029
rect 159477 160029 159493 160307
rect 159771 160029 159787 160307
rect 159477 142307 159787 160029
rect 159477 142029 159493 142307
rect 159771 142029 159787 142307
rect 159477 124307 159787 142029
rect 159477 124029 159493 124307
rect 159771 124029 159787 124307
rect 159477 106307 159787 124029
rect 159477 106029 159493 106307
rect 159771 106029 159787 106307
rect 159477 88307 159787 106029
rect 159477 88029 159493 88307
rect 159771 88029 159787 88307
rect 159477 70307 159787 88029
rect 159477 70029 159493 70307
rect 159771 70029 159787 70307
rect 159477 52307 159787 70029
rect 159477 52029 159493 52307
rect 159771 52029 159787 52307
rect 159477 34307 159787 52029
rect 159477 34029 159493 34307
rect 159771 34029 159787 34307
rect 159477 16307 159787 34029
rect 159477 16029 159493 16307
rect 159771 16029 159787 16307
rect 150477 -3331 150493 -3053
rect 150771 -3331 150787 -3053
rect 150477 -3827 150787 -3331
rect 159477 -3533 159787 16029
rect 162897 352419 163207 352915
rect 162897 352141 162913 352419
rect 163191 352141 163207 352419
rect 162897 343727 163207 352141
rect 162897 343449 162913 343727
rect 163191 343449 163207 343727
rect 162897 325727 163207 343449
rect 162897 325449 162913 325727
rect 163191 325449 163207 325727
rect 162897 307727 163207 325449
rect 162897 307449 162913 307727
rect 163191 307449 163207 307727
rect 162897 289727 163207 307449
rect 162897 289449 162913 289727
rect 163191 289449 163207 289727
rect 162897 271727 163207 289449
rect 162897 271449 162913 271727
rect 163191 271449 163207 271727
rect 162897 253727 163207 271449
rect 162897 253449 162913 253727
rect 163191 253449 163207 253727
rect 162897 235727 163207 253449
rect 162897 235449 162913 235727
rect 163191 235449 163207 235727
rect 162897 217727 163207 235449
rect 162897 217449 162913 217727
rect 163191 217449 163207 217727
rect 162897 199727 163207 217449
rect 162897 199449 162913 199727
rect 163191 199449 163207 199727
rect 162897 181727 163207 199449
rect 162897 181449 162913 181727
rect 163191 181449 163207 181727
rect 162897 163727 163207 181449
rect 162897 163449 162913 163727
rect 163191 163449 163207 163727
rect 162897 145727 163207 163449
rect 162897 145449 162913 145727
rect 163191 145449 163207 145727
rect 162897 127727 163207 145449
rect 162897 127449 162913 127727
rect 163191 127449 163207 127727
rect 162897 109727 163207 127449
rect 162897 109449 162913 109727
rect 163191 109449 163207 109727
rect 162897 91727 163207 109449
rect 162897 91449 162913 91727
rect 163191 91449 163207 91727
rect 162897 73727 163207 91449
rect 162897 73449 162913 73727
rect 163191 73449 163207 73727
rect 162897 55727 163207 73449
rect 162897 55449 162913 55727
rect 163191 55449 163207 55727
rect 162897 37727 163207 55449
rect 162897 37449 162913 37727
rect 163191 37449 163207 37727
rect 162897 19727 163207 37449
rect 162897 19449 162913 19727
rect 163191 19449 163207 19727
rect 162897 1727 163207 19449
rect 162897 1449 162913 1727
rect 163191 1449 163207 1727
rect 162897 -173 163207 1449
rect 162897 -451 162913 -173
rect 163191 -451 163207 -173
rect 162897 -947 163207 -451
rect 164757 345587 165067 353101
rect 164757 345309 164773 345587
rect 165051 345309 165067 345587
rect 164757 327587 165067 345309
rect 164757 327309 164773 327587
rect 165051 327309 165067 327587
rect 164757 309587 165067 327309
rect 164757 309309 164773 309587
rect 165051 309309 165067 309587
rect 164757 291587 165067 309309
rect 164757 291309 164773 291587
rect 165051 291309 165067 291587
rect 164757 273587 165067 291309
rect 164757 273309 164773 273587
rect 165051 273309 165067 273587
rect 164757 255587 165067 273309
rect 164757 255309 164773 255587
rect 165051 255309 165067 255587
rect 164757 237587 165067 255309
rect 164757 237309 164773 237587
rect 165051 237309 165067 237587
rect 164757 219587 165067 237309
rect 164757 219309 164773 219587
rect 165051 219309 165067 219587
rect 164757 201587 165067 219309
rect 164757 201309 164773 201587
rect 165051 201309 165067 201587
rect 164757 183587 165067 201309
rect 164757 183309 164773 183587
rect 165051 183309 165067 183587
rect 164757 165587 165067 183309
rect 164757 165309 164773 165587
rect 165051 165309 165067 165587
rect 164757 147587 165067 165309
rect 164757 147309 164773 147587
rect 165051 147309 165067 147587
rect 164757 129587 165067 147309
rect 164757 129309 164773 129587
rect 165051 129309 165067 129587
rect 164757 111587 165067 129309
rect 164757 111309 164773 111587
rect 165051 111309 165067 111587
rect 164757 93587 165067 111309
rect 164757 93309 164773 93587
rect 165051 93309 165067 93587
rect 164757 75587 165067 93309
rect 164757 75309 164773 75587
rect 165051 75309 165067 75587
rect 164757 57587 165067 75309
rect 164757 57309 164773 57587
rect 165051 57309 165067 57587
rect 164757 39587 165067 57309
rect 164757 39309 164773 39587
rect 165051 39309 165067 39587
rect 164757 21587 165067 39309
rect 164757 21309 164773 21587
rect 165051 21309 165067 21587
rect 164757 3587 165067 21309
rect 164757 3309 164773 3587
rect 165051 3309 165067 3587
rect 164757 -1133 165067 3309
rect 164757 -1411 164773 -1133
rect 165051 -1411 165067 -1133
rect 164757 -1907 165067 -1411
rect 166617 347447 166927 354061
rect 166617 347169 166633 347447
rect 166911 347169 166927 347447
rect 166617 329447 166927 347169
rect 166617 329169 166633 329447
rect 166911 329169 166927 329447
rect 166617 311447 166927 329169
rect 166617 311169 166633 311447
rect 166911 311169 166927 311447
rect 166617 293447 166927 311169
rect 166617 293169 166633 293447
rect 166911 293169 166927 293447
rect 166617 275447 166927 293169
rect 166617 275169 166633 275447
rect 166911 275169 166927 275447
rect 166617 257447 166927 275169
rect 166617 257169 166633 257447
rect 166911 257169 166927 257447
rect 166617 239447 166927 257169
rect 166617 239169 166633 239447
rect 166911 239169 166927 239447
rect 166617 221447 166927 239169
rect 166617 221169 166633 221447
rect 166911 221169 166927 221447
rect 166617 203447 166927 221169
rect 166617 203169 166633 203447
rect 166911 203169 166927 203447
rect 166617 185447 166927 203169
rect 166617 185169 166633 185447
rect 166911 185169 166927 185447
rect 166617 167447 166927 185169
rect 166617 167169 166633 167447
rect 166911 167169 166927 167447
rect 166617 149447 166927 167169
rect 166617 149169 166633 149447
rect 166911 149169 166927 149447
rect 166617 131447 166927 149169
rect 166617 131169 166633 131447
rect 166911 131169 166927 131447
rect 166617 113447 166927 131169
rect 166617 113169 166633 113447
rect 166911 113169 166927 113447
rect 166617 95447 166927 113169
rect 166617 95169 166633 95447
rect 166911 95169 166927 95447
rect 166617 77447 166927 95169
rect 166617 77169 166633 77447
rect 166911 77169 166927 77447
rect 166617 59447 166927 77169
rect 166617 59169 166633 59447
rect 166911 59169 166927 59447
rect 166617 41447 166927 59169
rect 166617 41169 166633 41447
rect 166911 41169 166927 41447
rect 166617 23447 166927 41169
rect 166617 23169 166633 23447
rect 166911 23169 166927 23447
rect 166617 5447 166927 23169
rect 166617 5169 166633 5447
rect 166911 5169 166927 5447
rect 166617 -2093 166927 5169
rect 166617 -2371 166633 -2093
rect 166911 -2371 166927 -2093
rect 166617 -2867 166927 -2371
rect 168477 349307 168787 355021
rect 177477 355779 177787 355795
rect 177477 355501 177493 355779
rect 177771 355501 177787 355779
rect 175617 354819 175927 354835
rect 175617 354541 175633 354819
rect 175911 354541 175927 354819
rect 173757 353859 174067 353875
rect 173757 353581 173773 353859
rect 174051 353581 174067 353859
rect 168477 349029 168493 349307
rect 168771 349029 168787 349307
rect 168477 331307 168787 349029
rect 168477 331029 168493 331307
rect 168771 331029 168787 331307
rect 168477 313307 168787 331029
rect 168477 313029 168493 313307
rect 168771 313029 168787 313307
rect 168477 295307 168787 313029
rect 168477 295029 168493 295307
rect 168771 295029 168787 295307
rect 168477 277307 168787 295029
rect 168477 277029 168493 277307
rect 168771 277029 168787 277307
rect 168477 259307 168787 277029
rect 168477 259029 168493 259307
rect 168771 259029 168787 259307
rect 168477 241307 168787 259029
rect 168477 241029 168493 241307
rect 168771 241029 168787 241307
rect 168477 223307 168787 241029
rect 168477 223029 168493 223307
rect 168771 223029 168787 223307
rect 168477 205307 168787 223029
rect 168477 205029 168493 205307
rect 168771 205029 168787 205307
rect 168477 187307 168787 205029
rect 168477 187029 168493 187307
rect 168771 187029 168787 187307
rect 168477 169307 168787 187029
rect 168477 169029 168493 169307
rect 168771 169029 168787 169307
rect 168477 151307 168787 169029
rect 168477 151029 168493 151307
rect 168771 151029 168787 151307
rect 168477 133307 168787 151029
rect 168477 133029 168493 133307
rect 168771 133029 168787 133307
rect 168477 115307 168787 133029
rect 168477 115029 168493 115307
rect 168771 115029 168787 115307
rect 168477 97307 168787 115029
rect 168477 97029 168493 97307
rect 168771 97029 168787 97307
rect 168477 79307 168787 97029
rect 168477 79029 168493 79307
rect 168771 79029 168787 79307
rect 168477 61307 168787 79029
rect 168477 61029 168493 61307
rect 168771 61029 168787 61307
rect 168477 43307 168787 61029
rect 168477 43029 168493 43307
rect 168771 43029 168787 43307
rect 168477 25307 168787 43029
rect 168477 25029 168493 25307
rect 168771 25029 168787 25307
rect 168477 7307 168787 25029
rect 168477 7029 168493 7307
rect 168771 7029 168787 7307
rect 159477 -3811 159493 -3533
rect 159771 -3811 159787 -3533
rect 159477 -3827 159787 -3811
rect 168477 -3053 168787 7029
rect 171897 352899 172207 352915
rect 171897 352621 171913 352899
rect 172191 352621 172207 352899
rect 171897 334727 172207 352621
rect 171897 334449 171913 334727
rect 172191 334449 172207 334727
rect 171897 316727 172207 334449
rect 171897 316449 171913 316727
rect 172191 316449 172207 316727
rect 171897 298727 172207 316449
rect 171897 298449 171913 298727
rect 172191 298449 172207 298727
rect 171897 280727 172207 298449
rect 171897 280449 171913 280727
rect 172191 280449 172207 280727
rect 171897 262727 172207 280449
rect 171897 262449 171913 262727
rect 172191 262449 172207 262727
rect 171897 244727 172207 262449
rect 171897 244449 171913 244727
rect 172191 244449 172207 244727
rect 171897 226727 172207 244449
rect 171897 226449 171913 226727
rect 172191 226449 172207 226727
rect 171897 208727 172207 226449
rect 171897 208449 171913 208727
rect 172191 208449 172207 208727
rect 171897 190727 172207 208449
rect 171897 190449 171913 190727
rect 172191 190449 172207 190727
rect 171897 172727 172207 190449
rect 171897 172449 171913 172727
rect 172191 172449 172207 172727
rect 171897 154727 172207 172449
rect 171897 154449 171913 154727
rect 172191 154449 172207 154727
rect 171897 136727 172207 154449
rect 171897 136449 171913 136727
rect 172191 136449 172207 136727
rect 171897 118727 172207 136449
rect 171897 118449 171913 118727
rect 172191 118449 172207 118727
rect 171897 100727 172207 118449
rect 171897 100449 171913 100727
rect 172191 100449 172207 100727
rect 171897 82727 172207 100449
rect 171897 82449 171913 82727
rect 172191 82449 172207 82727
rect 171897 64727 172207 82449
rect 171897 64449 171913 64727
rect 172191 64449 172207 64727
rect 171897 46727 172207 64449
rect 171897 46449 171913 46727
rect 172191 46449 172207 46727
rect 171897 28727 172207 46449
rect 171897 28449 171913 28727
rect 172191 28449 172207 28727
rect 171897 10727 172207 28449
rect 171897 10449 171913 10727
rect 172191 10449 172207 10727
rect 171897 -653 172207 10449
rect 171897 -931 171913 -653
rect 172191 -931 172207 -653
rect 171897 -947 172207 -931
rect 173757 336587 174067 353581
rect 173757 336309 173773 336587
rect 174051 336309 174067 336587
rect 173757 318587 174067 336309
rect 173757 318309 173773 318587
rect 174051 318309 174067 318587
rect 173757 300587 174067 318309
rect 173757 300309 173773 300587
rect 174051 300309 174067 300587
rect 173757 282587 174067 300309
rect 173757 282309 173773 282587
rect 174051 282309 174067 282587
rect 173757 264587 174067 282309
rect 173757 264309 173773 264587
rect 174051 264309 174067 264587
rect 173757 246587 174067 264309
rect 173757 246309 173773 246587
rect 174051 246309 174067 246587
rect 173757 228587 174067 246309
rect 173757 228309 173773 228587
rect 174051 228309 174067 228587
rect 173757 210587 174067 228309
rect 173757 210309 173773 210587
rect 174051 210309 174067 210587
rect 173757 192587 174067 210309
rect 173757 192309 173773 192587
rect 174051 192309 174067 192587
rect 173757 174587 174067 192309
rect 173757 174309 173773 174587
rect 174051 174309 174067 174587
rect 173757 156587 174067 174309
rect 173757 156309 173773 156587
rect 174051 156309 174067 156587
rect 173757 138587 174067 156309
rect 173757 138309 173773 138587
rect 174051 138309 174067 138587
rect 173757 120587 174067 138309
rect 173757 120309 173773 120587
rect 174051 120309 174067 120587
rect 173757 102587 174067 120309
rect 173757 102309 173773 102587
rect 174051 102309 174067 102587
rect 173757 84587 174067 102309
rect 173757 84309 173773 84587
rect 174051 84309 174067 84587
rect 173757 66587 174067 84309
rect 173757 66309 173773 66587
rect 174051 66309 174067 66587
rect 173757 48587 174067 66309
rect 173757 48309 173773 48587
rect 174051 48309 174067 48587
rect 173757 30587 174067 48309
rect 173757 30309 173773 30587
rect 174051 30309 174067 30587
rect 173757 12587 174067 30309
rect 173757 12309 173773 12587
rect 174051 12309 174067 12587
rect 173757 -1613 174067 12309
rect 173757 -1891 173773 -1613
rect 174051 -1891 174067 -1613
rect 173757 -1907 174067 -1891
rect 175617 338447 175927 354541
rect 175617 338169 175633 338447
rect 175911 338169 175927 338447
rect 175617 320447 175927 338169
rect 175617 320169 175633 320447
rect 175911 320169 175927 320447
rect 175617 302447 175927 320169
rect 175617 302169 175633 302447
rect 175911 302169 175927 302447
rect 175617 284447 175927 302169
rect 175617 284169 175633 284447
rect 175911 284169 175927 284447
rect 175617 266447 175927 284169
rect 175617 266169 175633 266447
rect 175911 266169 175927 266447
rect 175617 248447 175927 266169
rect 175617 248169 175633 248447
rect 175911 248169 175927 248447
rect 175617 230447 175927 248169
rect 175617 230169 175633 230447
rect 175911 230169 175927 230447
rect 175617 212447 175927 230169
rect 175617 212169 175633 212447
rect 175911 212169 175927 212447
rect 175617 194447 175927 212169
rect 175617 194169 175633 194447
rect 175911 194169 175927 194447
rect 175617 176447 175927 194169
rect 175617 176169 175633 176447
rect 175911 176169 175927 176447
rect 175617 158447 175927 176169
rect 175617 158169 175633 158447
rect 175911 158169 175927 158447
rect 175617 140447 175927 158169
rect 175617 140169 175633 140447
rect 175911 140169 175927 140447
rect 175617 122447 175927 140169
rect 175617 122169 175633 122447
rect 175911 122169 175927 122447
rect 175617 104447 175927 122169
rect 175617 104169 175633 104447
rect 175911 104169 175927 104447
rect 175617 86447 175927 104169
rect 175617 86169 175633 86447
rect 175911 86169 175927 86447
rect 175617 68447 175927 86169
rect 175617 68169 175633 68447
rect 175911 68169 175927 68447
rect 175617 50447 175927 68169
rect 175617 50169 175633 50447
rect 175911 50169 175927 50447
rect 175617 32447 175927 50169
rect 175617 32169 175633 32447
rect 175911 32169 175927 32447
rect 175617 14447 175927 32169
rect 175617 14169 175633 14447
rect 175911 14169 175927 14447
rect 175617 -2573 175927 14169
rect 175617 -2851 175633 -2573
rect 175911 -2851 175927 -2573
rect 175617 -2867 175927 -2851
rect 177477 340307 177787 355501
rect 186477 355299 186787 355795
rect 186477 355021 186493 355299
rect 186771 355021 186787 355299
rect 184617 354339 184927 354835
rect 184617 354061 184633 354339
rect 184911 354061 184927 354339
rect 182757 353379 183067 353875
rect 182757 353101 182773 353379
rect 183051 353101 183067 353379
rect 177477 340029 177493 340307
rect 177771 340029 177787 340307
rect 177477 322307 177787 340029
rect 177477 322029 177493 322307
rect 177771 322029 177787 322307
rect 177477 304307 177787 322029
rect 177477 304029 177493 304307
rect 177771 304029 177787 304307
rect 177477 286307 177787 304029
rect 177477 286029 177493 286307
rect 177771 286029 177787 286307
rect 177477 268307 177787 286029
rect 177477 268029 177493 268307
rect 177771 268029 177787 268307
rect 177477 250307 177787 268029
rect 177477 250029 177493 250307
rect 177771 250029 177787 250307
rect 177477 232307 177787 250029
rect 177477 232029 177493 232307
rect 177771 232029 177787 232307
rect 177477 214307 177787 232029
rect 177477 214029 177493 214307
rect 177771 214029 177787 214307
rect 177477 196307 177787 214029
rect 177477 196029 177493 196307
rect 177771 196029 177787 196307
rect 177477 178307 177787 196029
rect 177477 178029 177493 178307
rect 177771 178029 177787 178307
rect 177477 160307 177787 178029
rect 177477 160029 177493 160307
rect 177771 160029 177787 160307
rect 177477 142307 177787 160029
rect 177477 142029 177493 142307
rect 177771 142029 177787 142307
rect 177477 124307 177787 142029
rect 177477 124029 177493 124307
rect 177771 124029 177787 124307
rect 177477 106307 177787 124029
rect 177477 106029 177493 106307
rect 177771 106029 177787 106307
rect 177477 88307 177787 106029
rect 177477 88029 177493 88307
rect 177771 88029 177787 88307
rect 177477 70307 177787 88029
rect 177477 70029 177493 70307
rect 177771 70029 177787 70307
rect 177477 52307 177787 70029
rect 177477 52029 177493 52307
rect 177771 52029 177787 52307
rect 177477 34307 177787 52029
rect 177477 34029 177493 34307
rect 177771 34029 177787 34307
rect 177477 16307 177787 34029
rect 177477 16029 177493 16307
rect 177771 16029 177787 16307
rect 168477 -3331 168493 -3053
rect 168771 -3331 168787 -3053
rect 168477 -3827 168787 -3331
rect 177477 -3533 177787 16029
rect 180897 352419 181207 352915
rect 180897 352141 180913 352419
rect 181191 352141 181207 352419
rect 180897 343727 181207 352141
rect 180897 343449 180913 343727
rect 181191 343449 181207 343727
rect 180897 325727 181207 343449
rect 180897 325449 180913 325727
rect 181191 325449 181207 325727
rect 180897 307727 181207 325449
rect 180897 307449 180913 307727
rect 181191 307449 181207 307727
rect 180897 289727 181207 307449
rect 180897 289449 180913 289727
rect 181191 289449 181207 289727
rect 180897 271727 181207 289449
rect 180897 271449 180913 271727
rect 181191 271449 181207 271727
rect 180897 253727 181207 271449
rect 180897 253449 180913 253727
rect 181191 253449 181207 253727
rect 180897 235727 181207 253449
rect 180897 235449 180913 235727
rect 181191 235449 181207 235727
rect 180897 217727 181207 235449
rect 180897 217449 180913 217727
rect 181191 217449 181207 217727
rect 180897 199727 181207 217449
rect 180897 199449 180913 199727
rect 181191 199449 181207 199727
rect 180897 181727 181207 199449
rect 180897 181449 180913 181727
rect 181191 181449 181207 181727
rect 180897 163727 181207 181449
rect 180897 163449 180913 163727
rect 181191 163449 181207 163727
rect 180897 145727 181207 163449
rect 180897 145449 180913 145727
rect 181191 145449 181207 145727
rect 180897 127727 181207 145449
rect 180897 127449 180913 127727
rect 181191 127449 181207 127727
rect 180897 109727 181207 127449
rect 180897 109449 180913 109727
rect 181191 109449 181207 109727
rect 180897 91727 181207 109449
rect 180897 91449 180913 91727
rect 181191 91449 181207 91727
rect 180897 73727 181207 91449
rect 180897 73449 180913 73727
rect 181191 73449 181207 73727
rect 180897 55727 181207 73449
rect 180897 55449 180913 55727
rect 181191 55449 181207 55727
rect 180897 37727 181207 55449
rect 180897 37449 180913 37727
rect 181191 37449 181207 37727
rect 180897 19727 181207 37449
rect 180897 19449 180913 19727
rect 181191 19449 181207 19727
rect 180897 1727 181207 19449
rect 180897 1449 180913 1727
rect 181191 1449 181207 1727
rect 180897 -173 181207 1449
rect 180897 -451 180913 -173
rect 181191 -451 181207 -173
rect 180897 -947 181207 -451
rect 182757 345587 183067 353101
rect 182757 345309 182773 345587
rect 183051 345309 183067 345587
rect 182757 327587 183067 345309
rect 182757 327309 182773 327587
rect 183051 327309 183067 327587
rect 182757 309587 183067 327309
rect 182757 309309 182773 309587
rect 183051 309309 183067 309587
rect 182757 291587 183067 309309
rect 182757 291309 182773 291587
rect 183051 291309 183067 291587
rect 182757 273587 183067 291309
rect 182757 273309 182773 273587
rect 183051 273309 183067 273587
rect 182757 255587 183067 273309
rect 182757 255309 182773 255587
rect 183051 255309 183067 255587
rect 182757 237587 183067 255309
rect 182757 237309 182773 237587
rect 183051 237309 183067 237587
rect 182757 219587 183067 237309
rect 182757 219309 182773 219587
rect 183051 219309 183067 219587
rect 182757 201587 183067 219309
rect 182757 201309 182773 201587
rect 183051 201309 183067 201587
rect 182757 183587 183067 201309
rect 182757 183309 182773 183587
rect 183051 183309 183067 183587
rect 182757 165587 183067 183309
rect 182757 165309 182773 165587
rect 183051 165309 183067 165587
rect 182757 147587 183067 165309
rect 182757 147309 182773 147587
rect 183051 147309 183067 147587
rect 182757 129587 183067 147309
rect 182757 129309 182773 129587
rect 183051 129309 183067 129587
rect 182757 111587 183067 129309
rect 182757 111309 182773 111587
rect 183051 111309 183067 111587
rect 182757 93587 183067 111309
rect 182757 93309 182773 93587
rect 183051 93309 183067 93587
rect 182757 75587 183067 93309
rect 182757 75309 182773 75587
rect 183051 75309 183067 75587
rect 182757 57587 183067 75309
rect 182757 57309 182773 57587
rect 183051 57309 183067 57587
rect 182757 39587 183067 57309
rect 182757 39309 182773 39587
rect 183051 39309 183067 39587
rect 182757 21587 183067 39309
rect 182757 21309 182773 21587
rect 183051 21309 183067 21587
rect 182757 3587 183067 21309
rect 182757 3309 182773 3587
rect 183051 3309 183067 3587
rect 182757 -1133 183067 3309
rect 182757 -1411 182773 -1133
rect 183051 -1411 183067 -1133
rect 182757 -1907 183067 -1411
rect 184617 347447 184927 354061
rect 184617 347169 184633 347447
rect 184911 347169 184927 347447
rect 184617 329447 184927 347169
rect 184617 329169 184633 329447
rect 184911 329169 184927 329447
rect 184617 311447 184927 329169
rect 184617 311169 184633 311447
rect 184911 311169 184927 311447
rect 184617 293447 184927 311169
rect 184617 293169 184633 293447
rect 184911 293169 184927 293447
rect 184617 275447 184927 293169
rect 184617 275169 184633 275447
rect 184911 275169 184927 275447
rect 184617 257447 184927 275169
rect 184617 257169 184633 257447
rect 184911 257169 184927 257447
rect 184617 239447 184927 257169
rect 184617 239169 184633 239447
rect 184911 239169 184927 239447
rect 184617 221447 184927 239169
rect 184617 221169 184633 221447
rect 184911 221169 184927 221447
rect 184617 203447 184927 221169
rect 184617 203169 184633 203447
rect 184911 203169 184927 203447
rect 184617 185447 184927 203169
rect 184617 185169 184633 185447
rect 184911 185169 184927 185447
rect 184617 167447 184927 185169
rect 184617 167169 184633 167447
rect 184911 167169 184927 167447
rect 184617 149447 184927 167169
rect 184617 149169 184633 149447
rect 184911 149169 184927 149447
rect 184617 131447 184927 149169
rect 184617 131169 184633 131447
rect 184911 131169 184927 131447
rect 184617 113447 184927 131169
rect 184617 113169 184633 113447
rect 184911 113169 184927 113447
rect 184617 95447 184927 113169
rect 184617 95169 184633 95447
rect 184911 95169 184927 95447
rect 184617 77447 184927 95169
rect 184617 77169 184633 77447
rect 184911 77169 184927 77447
rect 184617 59447 184927 77169
rect 184617 59169 184633 59447
rect 184911 59169 184927 59447
rect 184617 41447 184927 59169
rect 184617 41169 184633 41447
rect 184911 41169 184927 41447
rect 184617 23447 184927 41169
rect 184617 23169 184633 23447
rect 184911 23169 184927 23447
rect 184617 5447 184927 23169
rect 184617 5169 184633 5447
rect 184911 5169 184927 5447
rect 184617 -2093 184927 5169
rect 184617 -2371 184633 -2093
rect 184911 -2371 184927 -2093
rect 184617 -2867 184927 -2371
rect 186477 349307 186787 355021
rect 195477 355779 195787 355795
rect 195477 355501 195493 355779
rect 195771 355501 195787 355779
rect 193617 354819 193927 354835
rect 193617 354541 193633 354819
rect 193911 354541 193927 354819
rect 191757 353859 192067 353875
rect 191757 353581 191773 353859
rect 192051 353581 192067 353859
rect 186477 349029 186493 349307
rect 186771 349029 186787 349307
rect 186477 331307 186787 349029
rect 186477 331029 186493 331307
rect 186771 331029 186787 331307
rect 186477 313307 186787 331029
rect 186477 313029 186493 313307
rect 186771 313029 186787 313307
rect 186477 295307 186787 313029
rect 186477 295029 186493 295307
rect 186771 295029 186787 295307
rect 186477 277307 186787 295029
rect 186477 277029 186493 277307
rect 186771 277029 186787 277307
rect 186477 259307 186787 277029
rect 186477 259029 186493 259307
rect 186771 259029 186787 259307
rect 186477 241307 186787 259029
rect 186477 241029 186493 241307
rect 186771 241029 186787 241307
rect 186477 223307 186787 241029
rect 186477 223029 186493 223307
rect 186771 223029 186787 223307
rect 186477 205307 186787 223029
rect 186477 205029 186493 205307
rect 186771 205029 186787 205307
rect 186477 187307 186787 205029
rect 186477 187029 186493 187307
rect 186771 187029 186787 187307
rect 186477 169307 186787 187029
rect 186477 169029 186493 169307
rect 186771 169029 186787 169307
rect 186477 151307 186787 169029
rect 186477 151029 186493 151307
rect 186771 151029 186787 151307
rect 186477 133307 186787 151029
rect 186477 133029 186493 133307
rect 186771 133029 186787 133307
rect 186477 115307 186787 133029
rect 186477 115029 186493 115307
rect 186771 115029 186787 115307
rect 186477 97307 186787 115029
rect 186477 97029 186493 97307
rect 186771 97029 186787 97307
rect 186477 79307 186787 97029
rect 186477 79029 186493 79307
rect 186771 79029 186787 79307
rect 186477 61307 186787 79029
rect 186477 61029 186493 61307
rect 186771 61029 186787 61307
rect 186477 43307 186787 61029
rect 186477 43029 186493 43307
rect 186771 43029 186787 43307
rect 186477 25307 186787 43029
rect 186477 25029 186493 25307
rect 186771 25029 186787 25307
rect 186477 7307 186787 25029
rect 186477 7029 186493 7307
rect 186771 7029 186787 7307
rect 177477 -3811 177493 -3533
rect 177771 -3811 177787 -3533
rect 177477 -3827 177787 -3811
rect 186477 -3053 186787 7029
rect 189897 352899 190207 352915
rect 189897 352621 189913 352899
rect 190191 352621 190207 352899
rect 189897 334727 190207 352621
rect 189897 334449 189913 334727
rect 190191 334449 190207 334727
rect 189897 316727 190207 334449
rect 189897 316449 189913 316727
rect 190191 316449 190207 316727
rect 189897 298727 190207 316449
rect 189897 298449 189913 298727
rect 190191 298449 190207 298727
rect 189897 280727 190207 298449
rect 189897 280449 189913 280727
rect 190191 280449 190207 280727
rect 189897 262727 190207 280449
rect 189897 262449 189913 262727
rect 190191 262449 190207 262727
rect 189897 244727 190207 262449
rect 189897 244449 189913 244727
rect 190191 244449 190207 244727
rect 189897 226727 190207 244449
rect 189897 226449 189913 226727
rect 190191 226449 190207 226727
rect 189897 208727 190207 226449
rect 189897 208449 189913 208727
rect 190191 208449 190207 208727
rect 189897 190727 190207 208449
rect 189897 190449 189913 190727
rect 190191 190449 190207 190727
rect 189897 172727 190207 190449
rect 189897 172449 189913 172727
rect 190191 172449 190207 172727
rect 189897 154727 190207 172449
rect 189897 154449 189913 154727
rect 190191 154449 190207 154727
rect 189897 136727 190207 154449
rect 189897 136449 189913 136727
rect 190191 136449 190207 136727
rect 189897 118727 190207 136449
rect 189897 118449 189913 118727
rect 190191 118449 190207 118727
rect 189897 100727 190207 118449
rect 189897 100449 189913 100727
rect 190191 100449 190207 100727
rect 189897 82727 190207 100449
rect 189897 82449 189913 82727
rect 190191 82449 190207 82727
rect 189897 64727 190207 82449
rect 189897 64449 189913 64727
rect 190191 64449 190207 64727
rect 189897 46727 190207 64449
rect 189897 46449 189913 46727
rect 190191 46449 190207 46727
rect 189897 28727 190207 46449
rect 189897 28449 189913 28727
rect 190191 28449 190207 28727
rect 189897 10727 190207 28449
rect 189897 10449 189913 10727
rect 190191 10449 190207 10727
rect 189897 -653 190207 10449
rect 189897 -931 189913 -653
rect 190191 -931 190207 -653
rect 189897 -947 190207 -931
rect 191757 336587 192067 353581
rect 191757 336309 191773 336587
rect 192051 336309 192067 336587
rect 191757 318587 192067 336309
rect 191757 318309 191773 318587
rect 192051 318309 192067 318587
rect 191757 300587 192067 318309
rect 191757 300309 191773 300587
rect 192051 300309 192067 300587
rect 191757 282587 192067 300309
rect 191757 282309 191773 282587
rect 192051 282309 192067 282587
rect 191757 264587 192067 282309
rect 191757 264309 191773 264587
rect 192051 264309 192067 264587
rect 191757 246587 192067 264309
rect 191757 246309 191773 246587
rect 192051 246309 192067 246587
rect 191757 228587 192067 246309
rect 191757 228309 191773 228587
rect 192051 228309 192067 228587
rect 191757 210587 192067 228309
rect 191757 210309 191773 210587
rect 192051 210309 192067 210587
rect 191757 192587 192067 210309
rect 191757 192309 191773 192587
rect 192051 192309 192067 192587
rect 191757 174587 192067 192309
rect 191757 174309 191773 174587
rect 192051 174309 192067 174587
rect 191757 156587 192067 174309
rect 191757 156309 191773 156587
rect 192051 156309 192067 156587
rect 191757 138587 192067 156309
rect 191757 138309 191773 138587
rect 192051 138309 192067 138587
rect 191757 120587 192067 138309
rect 191757 120309 191773 120587
rect 192051 120309 192067 120587
rect 191757 102587 192067 120309
rect 191757 102309 191773 102587
rect 192051 102309 192067 102587
rect 191757 84587 192067 102309
rect 191757 84309 191773 84587
rect 192051 84309 192067 84587
rect 191757 66587 192067 84309
rect 191757 66309 191773 66587
rect 192051 66309 192067 66587
rect 191757 48587 192067 66309
rect 191757 48309 191773 48587
rect 192051 48309 192067 48587
rect 191757 30587 192067 48309
rect 191757 30309 191773 30587
rect 192051 30309 192067 30587
rect 191757 12587 192067 30309
rect 191757 12309 191773 12587
rect 192051 12309 192067 12587
rect 191757 -1613 192067 12309
rect 191757 -1891 191773 -1613
rect 192051 -1891 192067 -1613
rect 191757 -1907 192067 -1891
rect 193617 338447 193927 354541
rect 193617 338169 193633 338447
rect 193911 338169 193927 338447
rect 193617 320447 193927 338169
rect 193617 320169 193633 320447
rect 193911 320169 193927 320447
rect 193617 302447 193927 320169
rect 193617 302169 193633 302447
rect 193911 302169 193927 302447
rect 193617 284447 193927 302169
rect 193617 284169 193633 284447
rect 193911 284169 193927 284447
rect 193617 266447 193927 284169
rect 193617 266169 193633 266447
rect 193911 266169 193927 266447
rect 193617 248447 193927 266169
rect 193617 248169 193633 248447
rect 193911 248169 193927 248447
rect 193617 230447 193927 248169
rect 193617 230169 193633 230447
rect 193911 230169 193927 230447
rect 193617 212447 193927 230169
rect 193617 212169 193633 212447
rect 193911 212169 193927 212447
rect 193617 194447 193927 212169
rect 193617 194169 193633 194447
rect 193911 194169 193927 194447
rect 193617 176447 193927 194169
rect 193617 176169 193633 176447
rect 193911 176169 193927 176447
rect 193617 158447 193927 176169
rect 193617 158169 193633 158447
rect 193911 158169 193927 158447
rect 193617 140447 193927 158169
rect 193617 140169 193633 140447
rect 193911 140169 193927 140447
rect 193617 122447 193927 140169
rect 193617 122169 193633 122447
rect 193911 122169 193927 122447
rect 193617 104447 193927 122169
rect 193617 104169 193633 104447
rect 193911 104169 193927 104447
rect 193617 86447 193927 104169
rect 193617 86169 193633 86447
rect 193911 86169 193927 86447
rect 193617 68447 193927 86169
rect 193617 68169 193633 68447
rect 193911 68169 193927 68447
rect 193617 50447 193927 68169
rect 193617 50169 193633 50447
rect 193911 50169 193927 50447
rect 193617 32447 193927 50169
rect 193617 32169 193633 32447
rect 193911 32169 193927 32447
rect 193617 14447 193927 32169
rect 193617 14169 193633 14447
rect 193911 14169 193927 14447
rect 193617 -2573 193927 14169
rect 193617 -2851 193633 -2573
rect 193911 -2851 193927 -2573
rect 193617 -2867 193927 -2851
rect 195477 340307 195787 355501
rect 204477 355299 204787 355795
rect 204477 355021 204493 355299
rect 204771 355021 204787 355299
rect 202617 354339 202927 354835
rect 202617 354061 202633 354339
rect 202911 354061 202927 354339
rect 200757 353379 201067 353875
rect 200757 353101 200773 353379
rect 201051 353101 201067 353379
rect 195477 340029 195493 340307
rect 195771 340029 195787 340307
rect 195477 322307 195787 340029
rect 195477 322029 195493 322307
rect 195771 322029 195787 322307
rect 195477 304307 195787 322029
rect 195477 304029 195493 304307
rect 195771 304029 195787 304307
rect 195477 286307 195787 304029
rect 195477 286029 195493 286307
rect 195771 286029 195787 286307
rect 195477 268307 195787 286029
rect 195477 268029 195493 268307
rect 195771 268029 195787 268307
rect 195477 250307 195787 268029
rect 195477 250029 195493 250307
rect 195771 250029 195787 250307
rect 195477 232307 195787 250029
rect 195477 232029 195493 232307
rect 195771 232029 195787 232307
rect 195477 214307 195787 232029
rect 195477 214029 195493 214307
rect 195771 214029 195787 214307
rect 195477 196307 195787 214029
rect 195477 196029 195493 196307
rect 195771 196029 195787 196307
rect 195477 178307 195787 196029
rect 195477 178029 195493 178307
rect 195771 178029 195787 178307
rect 195477 160307 195787 178029
rect 195477 160029 195493 160307
rect 195771 160029 195787 160307
rect 195477 142307 195787 160029
rect 195477 142029 195493 142307
rect 195771 142029 195787 142307
rect 195477 124307 195787 142029
rect 195477 124029 195493 124307
rect 195771 124029 195787 124307
rect 195477 106307 195787 124029
rect 195477 106029 195493 106307
rect 195771 106029 195787 106307
rect 195477 88307 195787 106029
rect 195477 88029 195493 88307
rect 195771 88029 195787 88307
rect 195477 70307 195787 88029
rect 195477 70029 195493 70307
rect 195771 70029 195787 70307
rect 195477 52307 195787 70029
rect 195477 52029 195493 52307
rect 195771 52029 195787 52307
rect 195477 34307 195787 52029
rect 195477 34029 195493 34307
rect 195771 34029 195787 34307
rect 195477 16307 195787 34029
rect 195477 16029 195493 16307
rect 195771 16029 195787 16307
rect 186477 -3331 186493 -3053
rect 186771 -3331 186787 -3053
rect 186477 -3827 186787 -3331
rect 195477 -3533 195787 16029
rect 198897 352419 199207 352915
rect 198897 352141 198913 352419
rect 199191 352141 199207 352419
rect 198897 343727 199207 352141
rect 198897 343449 198913 343727
rect 199191 343449 199207 343727
rect 198897 325727 199207 343449
rect 198897 325449 198913 325727
rect 199191 325449 199207 325727
rect 198897 307727 199207 325449
rect 198897 307449 198913 307727
rect 199191 307449 199207 307727
rect 198897 289727 199207 307449
rect 198897 289449 198913 289727
rect 199191 289449 199207 289727
rect 198897 271727 199207 289449
rect 198897 271449 198913 271727
rect 199191 271449 199207 271727
rect 198897 253727 199207 271449
rect 198897 253449 198913 253727
rect 199191 253449 199207 253727
rect 198897 235727 199207 253449
rect 198897 235449 198913 235727
rect 199191 235449 199207 235727
rect 198897 217727 199207 235449
rect 198897 217449 198913 217727
rect 199191 217449 199207 217727
rect 198897 199727 199207 217449
rect 198897 199449 198913 199727
rect 199191 199449 199207 199727
rect 198897 181727 199207 199449
rect 198897 181449 198913 181727
rect 199191 181449 199207 181727
rect 198897 163727 199207 181449
rect 198897 163449 198913 163727
rect 199191 163449 199207 163727
rect 198897 145727 199207 163449
rect 198897 145449 198913 145727
rect 199191 145449 199207 145727
rect 198897 127727 199207 145449
rect 198897 127449 198913 127727
rect 199191 127449 199207 127727
rect 198897 109727 199207 127449
rect 198897 109449 198913 109727
rect 199191 109449 199207 109727
rect 198897 91727 199207 109449
rect 198897 91449 198913 91727
rect 199191 91449 199207 91727
rect 198897 73727 199207 91449
rect 198897 73449 198913 73727
rect 199191 73449 199207 73727
rect 198897 55727 199207 73449
rect 198897 55449 198913 55727
rect 199191 55449 199207 55727
rect 198897 37727 199207 55449
rect 198897 37449 198913 37727
rect 199191 37449 199207 37727
rect 198897 19727 199207 37449
rect 198897 19449 198913 19727
rect 199191 19449 199207 19727
rect 198897 1727 199207 19449
rect 198897 1449 198913 1727
rect 199191 1449 199207 1727
rect 198897 -173 199207 1449
rect 198897 -451 198913 -173
rect 199191 -451 199207 -173
rect 198897 -947 199207 -451
rect 200757 345587 201067 353101
rect 200757 345309 200773 345587
rect 201051 345309 201067 345587
rect 200757 327587 201067 345309
rect 200757 327309 200773 327587
rect 201051 327309 201067 327587
rect 200757 309587 201067 327309
rect 200757 309309 200773 309587
rect 201051 309309 201067 309587
rect 200757 291587 201067 309309
rect 200757 291309 200773 291587
rect 201051 291309 201067 291587
rect 200757 273587 201067 291309
rect 200757 273309 200773 273587
rect 201051 273309 201067 273587
rect 200757 255587 201067 273309
rect 200757 255309 200773 255587
rect 201051 255309 201067 255587
rect 200757 237587 201067 255309
rect 200757 237309 200773 237587
rect 201051 237309 201067 237587
rect 200757 219587 201067 237309
rect 200757 219309 200773 219587
rect 201051 219309 201067 219587
rect 200757 201587 201067 219309
rect 200757 201309 200773 201587
rect 201051 201309 201067 201587
rect 200757 183587 201067 201309
rect 200757 183309 200773 183587
rect 201051 183309 201067 183587
rect 200757 165587 201067 183309
rect 200757 165309 200773 165587
rect 201051 165309 201067 165587
rect 200757 147587 201067 165309
rect 200757 147309 200773 147587
rect 201051 147309 201067 147587
rect 200757 129587 201067 147309
rect 200757 129309 200773 129587
rect 201051 129309 201067 129587
rect 200757 111587 201067 129309
rect 200757 111309 200773 111587
rect 201051 111309 201067 111587
rect 200757 93587 201067 111309
rect 200757 93309 200773 93587
rect 201051 93309 201067 93587
rect 200757 75587 201067 93309
rect 200757 75309 200773 75587
rect 201051 75309 201067 75587
rect 200757 57587 201067 75309
rect 200757 57309 200773 57587
rect 201051 57309 201067 57587
rect 200757 39587 201067 57309
rect 200757 39309 200773 39587
rect 201051 39309 201067 39587
rect 200757 21587 201067 39309
rect 200757 21309 200773 21587
rect 201051 21309 201067 21587
rect 200757 3587 201067 21309
rect 200757 3309 200773 3587
rect 201051 3309 201067 3587
rect 200757 -1133 201067 3309
rect 200757 -1411 200773 -1133
rect 201051 -1411 201067 -1133
rect 200757 -1907 201067 -1411
rect 202617 347447 202927 354061
rect 202617 347169 202633 347447
rect 202911 347169 202927 347447
rect 202617 329447 202927 347169
rect 202617 329169 202633 329447
rect 202911 329169 202927 329447
rect 202617 311447 202927 329169
rect 202617 311169 202633 311447
rect 202911 311169 202927 311447
rect 202617 293447 202927 311169
rect 202617 293169 202633 293447
rect 202911 293169 202927 293447
rect 202617 275447 202927 293169
rect 202617 275169 202633 275447
rect 202911 275169 202927 275447
rect 202617 257447 202927 275169
rect 202617 257169 202633 257447
rect 202911 257169 202927 257447
rect 202617 239447 202927 257169
rect 202617 239169 202633 239447
rect 202911 239169 202927 239447
rect 202617 221447 202927 239169
rect 202617 221169 202633 221447
rect 202911 221169 202927 221447
rect 202617 203447 202927 221169
rect 202617 203169 202633 203447
rect 202911 203169 202927 203447
rect 202617 185447 202927 203169
rect 202617 185169 202633 185447
rect 202911 185169 202927 185447
rect 202617 167447 202927 185169
rect 202617 167169 202633 167447
rect 202911 167169 202927 167447
rect 202617 149447 202927 167169
rect 202617 149169 202633 149447
rect 202911 149169 202927 149447
rect 202617 131447 202927 149169
rect 202617 131169 202633 131447
rect 202911 131169 202927 131447
rect 202617 113447 202927 131169
rect 202617 113169 202633 113447
rect 202911 113169 202927 113447
rect 202617 95447 202927 113169
rect 202617 95169 202633 95447
rect 202911 95169 202927 95447
rect 202617 77447 202927 95169
rect 202617 77169 202633 77447
rect 202911 77169 202927 77447
rect 202617 59447 202927 77169
rect 202617 59169 202633 59447
rect 202911 59169 202927 59447
rect 202617 41447 202927 59169
rect 202617 41169 202633 41447
rect 202911 41169 202927 41447
rect 202617 23447 202927 41169
rect 202617 23169 202633 23447
rect 202911 23169 202927 23447
rect 202617 5447 202927 23169
rect 202617 5169 202633 5447
rect 202911 5169 202927 5447
rect 202617 -2093 202927 5169
rect 202617 -2371 202633 -2093
rect 202911 -2371 202927 -2093
rect 202617 -2867 202927 -2371
rect 204477 349307 204787 355021
rect 213477 355779 213787 355795
rect 213477 355501 213493 355779
rect 213771 355501 213787 355779
rect 211617 354819 211927 354835
rect 211617 354541 211633 354819
rect 211911 354541 211927 354819
rect 209757 353859 210067 353875
rect 209757 353581 209773 353859
rect 210051 353581 210067 353859
rect 204477 349029 204493 349307
rect 204771 349029 204787 349307
rect 204477 331307 204787 349029
rect 204477 331029 204493 331307
rect 204771 331029 204787 331307
rect 204477 313307 204787 331029
rect 204477 313029 204493 313307
rect 204771 313029 204787 313307
rect 204477 295307 204787 313029
rect 204477 295029 204493 295307
rect 204771 295029 204787 295307
rect 204477 277307 204787 295029
rect 204477 277029 204493 277307
rect 204771 277029 204787 277307
rect 204477 259307 204787 277029
rect 204477 259029 204493 259307
rect 204771 259029 204787 259307
rect 204477 241307 204787 259029
rect 204477 241029 204493 241307
rect 204771 241029 204787 241307
rect 204477 223307 204787 241029
rect 204477 223029 204493 223307
rect 204771 223029 204787 223307
rect 204477 205307 204787 223029
rect 204477 205029 204493 205307
rect 204771 205029 204787 205307
rect 204477 187307 204787 205029
rect 204477 187029 204493 187307
rect 204771 187029 204787 187307
rect 204477 169307 204787 187029
rect 204477 169029 204493 169307
rect 204771 169029 204787 169307
rect 204477 151307 204787 169029
rect 204477 151029 204493 151307
rect 204771 151029 204787 151307
rect 204477 133307 204787 151029
rect 204477 133029 204493 133307
rect 204771 133029 204787 133307
rect 204477 115307 204787 133029
rect 204477 115029 204493 115307
rect 204771 115029 204787 115307
rect 204477 97307 204787 115029
rect 204477 97029 204493 97307
rect 204771 97029 204787 97307
rect 204477 79307 204787 97029
rect 204477 79029 204493 79307
rect 204771 79029 204787 79307
rect 204477 61307 204787 79029
rect 204477 61029 204493 61307
rect 204771 61029 204787 61307
rect 204477 43307 204787 61029
rect 204477 43029 204493 43307
rect 204771 43029 204787 43307
rect 204477 25307 204787 43029
rect 204477 25029 204493 25307
rect 204771 25029 204787 25307
rect 204477 7307 204787 25029
rect 204477 7029 204493 7307
rect 204771 7029 204787 7307
rect 195477 -3811 195493 -3533
rect 195771 -3811 195787 -3533
rect 195477 -3827 195787 -3811
rect 204477 -3053 204787 7029
rect 207897 352899 208207 352915
rect 207897 352621 207913 352899
rect 208191 352621 208207 352899
rect 207897 334727 208207 352621
rect 207897 334449 207913 334727
rect 208191 334449 208207 334727
rect 207897 316727 208207 334449
rect 207897 316449 207913 316727
rect 208191 316449 208207 316727
rect 207897 298727 208207 316449
rect 207897 298449 207913 298727
rect 208191 298449 208207 298727
rect 207897 280727 208207 298449
rect 207897 280449 207913 280727
rect 208191 280449 208207 280727
rect 207897 262727 208207 280449
rect 207897 262449 207913 262727
rect 208191 262449 208207 262727
rect 207897 244727 208207 262449
rect 207897 244449 207913 244727
rect 208191 244449 208207 244727
rect 207897 226727 208207 244449
rect 207897 226449 207913 226727
rect 208191 226449 208207 226727
rect 207897 208727 208207 226449
rect 207897 208449 207913 208727
rect 208191 208449 208207 208727
rect 207897 190727 208207 208449
rect 207897 190449 207913 190727
rect 208191 190449 208207 190727
rect 207897 172727 208207 190449
rect 207897 172449 207913 172727
rect 208191 172449 208207 172727
rect 207897 154727 208207 172449
rect 207897 154449 207913 154727
rect 208191 154449 208207 154727
rect 207897 136727 208207 154449
rect 207897 136449 207913 136727
rect 208191 136449 208207 136727
rect 207897 118727 208207 136449
rect 207897 118449 207913 118727
rect 208191 118449 208207 118727
rect 207897 100727 208207 118449
rect 207897 100449 207913 100727
rect 208191 100449 208207 100727
rect 207897 82727 208207 100449
rect 207897 82449 207913 82727
rect 208191 82449 208207 82727
rect 207897 64727 208207 82449
rect 207897 64449 207913 64727
rect 208191 64449 208207 64727
rect 207897 46727 208207 64449
rect 207897 46449 207913 46727
rect 208191 46449 208207 46727
rect 207897 28727 208207 46449
rect 207897 28449 207913 28727
rect 208191 28449 208207 28727
rect 207897 10727 208207 28449
rect 207897 10449 207913 10727
rect 208191 10449 208207 10727
rect 207897 -653 208207 10449
rect 207897 -931 207913 -653
rect 208191 -931 208207 -653
rect 207897 -947 208207 -931
rect 209757 336587 210067 353581
rect 209757 336309 209773 336587
rect 210051 336309 210067 336587
rect 209757 318587 210067 336309
rect 209757 318309 209773 318587
rect 210051 318309 210067 318587
rect 209757 300587 210067 318309
rect 209757 300309 209773 300587
rect 210051 300309 210067 300587
rect 209757 282587 210067 300309
rect 209757 282309 209773 282587
rect 210051 282309 210067 282587
rect 209757 264587 210067 282309
rect 209757 264309 209773 264587
rect 210051 264309 210067 264587
rect 209757 246587 210067 264309
rect 209757 246309 209773 246587
rect 210051 246309 210067 246587
rect 209757 228587 210067 246309
rect 209757 228309 209773 228587
rect 210051 228309 210067 228587
rect 209757 210587 210067 228309
rect 209757 210309 209773 210587
rect 210051 210309 210067 210587
rect 209757 192587 210067 210309
rect 209757 192309 209773 192587
rect 210051 192309 210067 192587
rect 209757 174587 210067 192309
rect 209757 174309 209773 174587
rect 210051 174309 210067 174587
rect 209757 156587 210067 174309
rect 209757 156309 209773 156587
rect 210051 156309 210067 156587
rect 209757 138587 210067 156309
rect 209757 138309 209773 138587
rect 210051 138309 210067 138587
rect 209757 120587 210067 138309
rect 209757 120309 209773 120587
rect 210051 120309 210067 120587
rect 209757 102587 210067 120309
rect 209757 102309 209773 102587
rect 210051 102309 210067 102587
rect 209757 84587 210067 102309
rect 209757 84309 209773 84587
rect 210051 84309 210067 84587
rect 209757 66587 210067 84309
rect 209757 66309 209773 66587
rect 210051 66309 210067 66587
rect 209757 48587 210067 66309
rect 209757 48309 209773 48587
rect 210051 48309 210067 48587
rect 209757 30587 210067 48309
rect 209757 30309 209773 30587
rect 210051 30309 210067 30587
rect 209757 12587 210067 30309
rect 209757 12309 209773 12587
rect 210051 12309 210067 12587
rect 209757 -1613 210067 12309
rect 209757 -1891 209773 -1613
rect 210051 -1891 210067 -1613
rect 209757 -1907 210067 -1891
rect 211617 338447 211927 354541
rect 211617 338169 211633 338447
rect 211911 338169 211927 338447
rect 211617 320447 211927 338169
rect 211617 320169 211633 320447
rect 211911 320169 211927 320447
rect 211617 302447 211927 320169
rect 211617 302169 211633 302447
rect 211911 302169 211927 302447
rect 211617 284447 211927 302169
rect 211617 284169 211633 284447
rect 211911 284169 211927 284447
rect 211617 266447 211927 284169
rect 211617 266169 211633 266447
rect 211911 266169 211927 266447
rect 211617 248447 211927 266169
rect 211617 248169 211633 248447
rect 211911 248169 211927 248447
rect 211617 230447 211927 248169
rect 211617 230169 211633 230447
rect 211911 230169 211927 230447
rect 211617 212447 211927 230169
rect 211617 212169 211633 212447
rect 211911 212169 211927 212447
rect 211617 194447 211927 212169
rect 211617 194169 211633 194447
rect 211911 194169 211927 194447
rect 211617 176447 211927 194169
rect 211617 176169 211633 176447
rect 211911 176169 211927 176447
rect 211617 158447 211927 176169
rect 211617 158169 211633 158447
rect 211911 158169 211927 158447
rect 211617 140447 211927 158169
rect 211617 140169 211633 140447
rect 211911 140169 211927 140447
rect 211617 122447 211927 140169
rect 211617 122169 211633 122447
rect 211911 122169 211927 122447
rect 211617 104447 211927 122169
rect 211617 104169 211633 104447
rect 211911 104169 211927 104447
rect 211617 86447 211927 104169
rect 211617 86169 211633 86447
rect 211911 86169 211927 86447
rect 211617 68447 211927 86169
rect 211617 68169 211633 68447
rect 211911 68169 211927 68447
rect 211617 50447 211927 68169
rect 211617 50169 211633 50447
rect 211911 50169 211927 50447
rect 211617 32447 211927 50169
rect 211617 32169 211633 32447
rect 211911 32169 211927 32447
rect 211617 14447 211927 32169
rect 211617 14169 211633 14447
rect 211911 14169 211927 14447
rect 211617 -2573 211927 14169
rect 211617 -2851 211633 -2573
rect 211911 -2851 211927 -2573
rect 211617 -2867 211927 -2851
rect 213477 340307 213787 355501
rect 222477 355299 222787 355795
rect 222477 355021 222493 355299
rect 222771 355021 222787 355299
rect 220617 354339 220927 354835
rect 220617 354061 220633 354339
rect 220911 354061 220927 354339
rect 218757 353379 219067 353875
rect 218757 353101 218773 353379
rect 219051 353101 219067 353379
rect 213477 340029 213493 340307
rect 213771 340029 213787 340307
rect 213477 322307 213787 340029
rect 213477 322029 213493 322307
rect 213771 322029 213787 322307
rect 213477 304307 213787 322029
rect 213477 304029 213493 304307
rect 213771 304029 213787 304307
rect 213477 286307 213787 304029
rect 213477 286029 213493 286307
rect 213771 286029 213787 286307
rect 213477 268307 213787 286029
rect 213477 268029 213493 268307
rect 213771 268029 213787 268307
rect 213477 250307 213787 268029
rect 213477 250029 213493 250307
rect 213771 250029 213787 250307
rect 213477 232307 213787 250029
rect 213477 232029 213493 232307
rect 213771 232029 213787 232307
rect 213477 214307 213787 232029
rect 213477 214029 213493 214307
rect 213771 214029 213787 214307
rect 213477 196307 213787 214029
rect 213477 196029 213493 196307
rect 213771 196029 213787 196307
rect 213477 178307 213787 196029
rect 213477 178029 213493 178307
rect 213771 178029 213787 178307
rect 213477 160307 213787 178029
rect 213477 160029 213493 160307
rect 213771 160029 213787 160307
rect 213477 142307 213787 160029
rect 213477 142029 213493 142307
rect 213771 142029 213787 142307
rect 213477 124307 213787 142029
rect 213477 124029 213493 124307
rect 213771 124029 213787 124307
rect 213477 106307 213787 124029
rect 213477 106029 213493 106307
rect 213771 106029 213787 106307
rect 213477 88307 213787 106029
rect 213477 88029 213493 88307
rect 213771 88029 213787 88307
rect 213477 70307 213787 88029
rect 213477 70029 213493 70307
rect 213771 70029 213787 70307
rect 213477 52307 213787 70029
rect 213477 52029 213493 52307
rect 213771 52029 213787 52307
rect 213477 34307 213787 52029
rect 213477 34029 213493 34307
rect 213771 34029 213787 34307
rect 213477 16307 213787 34029
rect 213477 16029 213493 16307
rect 213771 16029 213787 16307
rect 204477 -3331 204493 -3053
rect 204771 -3331 204787 -3053
rect 204477 -3827 204787 -3331
rect 213477 -3533 213787 16029
rect 216897 352419 217207 352915
rect 216897 352141 216913 352419
rect 217191 352141 217207 352419
rect 216897 343727 217207 352141
rect 216897 343449 216913 343727
rect 217191 343449 217207 343727
rect 216897 325727 217207 343449
rect 216897 325449 216913 325727
rect 217191 325449 217207 325727
rect 216897 307727 217207 325449
rect 216897 307449 216913 307727
rect 217191 307449 217207 307727
rect 216897 289727 217207 307449
rect 216897 289449 216913 289727
rect 217191 289449 217207 289727
rect 216897 271727 217207 289449
rect 216897 271449 216913 271727
rect 217191 271449 217207 271727
rect 216897 253727 217207 271449
rect 216897 253449 216913 253727
rect 217191 253449 217207 253727
rect 216897 235727 217207 253449
rect 216897 235449 216913 235727
rect 217191 235449 217207 235727
rect 216897 217727 217207 235449
rect 216897 217449 216913 217727
rect 217191 217449 217207 217727
rect 216897 199727 217207 217449
rect 216897 199449 216913 199727
rect 217191 199449 217207 199727
rect 216897 181727 217207 199449
rect 216897 181449 216913 181727
rect 217191 181449 217207 181727
rect 216897 163727 217207 181449
rect 216897 163449 216913 163727
rect 217191 163449 217207 163727
rect 216897 145727 217207 163449
rect 216897 145449 216913 145727
rect 217191 145449 217207 145727
rect 216897 127727 217207 145449
rect 216897 127449 216913 127727
rect 217191 127449 217207 127727
rect 216897 109727 217207 127449
rect 216897 109449 216913 109727
rect 217191 109449 217207 109727
rect 216897 91727 217207 109449
rect 216897 91449 216913 91727
rect 217191 91449 217207 91727
rect 216897 73727 217207 91449
rect 216897 73449 216913 73727
rect 217191 73449 217207 73727
rect 216897 55727 217207 73449
rect 216897 55449 216913 55727
rect 217191 55449 217207 55727
rect 216897 37727 217207 55449
rect 216897 37449 216913 37727
rect 217191 37449 217207 37727
rect 216897 19727 217207 37449
rect 216897 19449 216913 19727
rect 217191 19449 217207 19727
rect 216897 1727 217207 19449
rect 216897 1449 216913 1727
rect 217191 1449 217207 1727
rect 216897 -173 217207 1449
rect 216897 -451 216913 -173
rect 217191 -451 217207 -173
rect 216897 -947 217207 -451
rect 218757 345587 219067 353101
rect 218757 345309 218773 345587
rect 219051 345309 219067 345587
rect 218757 327587 219067 345309
rect 218757 327309 218773 327587
rect 219051 327309 219067 327587
rect 218757 309587 219067 327309
rect 218757 309309 218773 309587
rect 219051 309309 219067 309587
rect 218757 291587 219067 309309
rect 218757 291309 218773 291587
rect 219051 291309 219067 291587
rect 218757 273587 219067 291309
rect 218757 273309 218773 273587
rect 219051 273309 219067 273587
rect 218757 255587 219067 273309
rect 218757 255309 218773 255587
rect 219051 255309 219067 255587
rect 218757 237587 219067 255309
rect 218757 237309 218773 237587
rect 219051 237309 219067 237587
rect 218757 219587 219067 237309
rect 218757 219309 218773 219587
rect 219051 219309 219067 219587
rect 218757 201587 219067 219309
rect 218757 201309 218773 201587
rect 219051 201309 219067 201587
rect 218757 183587 219067 201309
rect 218757 183309 218773 183587
rect 219051 183309 219067 183587
rect 218757 165587 219067 183309
rect 218757 165309 218773 165587
rect 219051 165309 219067 165587
rect 218757 147587 219067 165309
rect 218757 147309 218773 147587
rect 219051 147309 219067 147587
rect 218757 129587 219067 147309
rect 218757 129309 218773 129587
rect 219051 129309 219067 129587
rect 218757 111587 219067 129309
rect 218757 111309 218773 111587
rect 219051 111309 219067 111587
rect 218757 93587 219067 111309
rect 218757 93309 218773 93587
rect 219051 93309 219067 93587
rect 218757 75587 219067 93309
rect 218757 75309 218773 75587
rect 219051 75309 219067 75587
rect 218757 57587 219067 75309
rect 218757 57309 218773 57587
rect 219051 57309 219067 57587
rect 218757 39587 219067 57309
rect 218757 39309 218773 39587
rect 219051 39309 219067 39587
rect 218757 21587 219067 39309
rect 218757 21309 218773 21587
rect 219051 21309 219067 21587
rect 218757 3587 219067 21309
rect 218757 3309 218773 3587
rect 219051 3309 219067 3587
rect 218757 -1133 219067 3309
rect 218757 -1411 218773 -1133
rect 219051 -1411 219067 -1133
rect 218757 -1907 219067 -1411
rect 220617 347447 220927 354061
rect 220617 347169 220633 347447
rect 220911 347169 220927 347447
rect 220617 329447 220927 347169
rect 220617 329169 220633 329447
rect 220911 329169 220927 329447
rect 220617 311447 220927 329169
rect 220617 311169 220633 311447
rect 220911 311169 220927 311447
rect 220617 293447 220927 311169
rect 220617 293169 220633 293447
rect 220911 293169 220927 293447
rect 220617 275447 220927 293169
rect 220617 275169 220633 275447
rect 220911 275169 220927 275447
rect 220617 257447 220927 275169
rect 220617 257169 220633 257447
rect 220911 257169 220927 257447
rect 220617 239447 220927 257169
rect 220617 239169 220633 239447
rect 220911 239169 220927 239447
rect 220617 221447 220927 239169
rect 220617 221169 220633 221447
rect 220911 221169 220927 221447
rect 220617 203447 220927 221169
rect 220617 203169 220633 203447
rect 220911 203169 220927 203447
rect 220617 185447 220927 203169
rect 220617 185169 220633 185447
rect 220911 185169 220927 185447
rect 220617 167447 220927 185169
rect 220617 167169 220633 167447
rect 220911 167169 220927 167447
rect 220617 149447 220927 167169
rect 220617 149169 220633 149447
rect 220911 149169 220927 149447
rect 220617 131447 220927 149169
rect 220617 131169 220633 131447
rect 220911 131169 220927 131447
rect 220617 113447 220927 131169
rect 220617 113169 220633 113447
rect 220911 113169 220927 113447
rect 220617 95447 220927 113169
rect 220617 95169 220633 95447
rect 220911 95169 220927 95447
rect 220617 77447 220927 95169
rect 220617 77169 220633 77447
rect 220911 77169 220927 77447
rect 220617 59447 220927 77169
rect 220617 59169 220633 59447
rect 220911 59169 220927 59447
rect 220617 41447 220927 59169
rect 220617 41169 220633 41447
rect 220911 41169 220927 41447
rect 220617 23447 220927 41169
rect 220617 23169 220633 23447
rect 220911 23169 220927 23447
rect 220617 5447 220927 23169
rect 220617 5169 220633 5447
rect 220911 5169 220927 5447
rect 220617 -2093 220927 5169
rect 220617 -2371 220633 -2093
rect 220911 -2371 220927 -2093
rect 220617 -2867 220927 -2371
rect 222477 349307 222787 355021
rect 231477 355779 231787 355795
rect 231477 355501 231493 355779
rect 231771 355501 231787 355779
rect 229617 354819 229927 354835
rect 229617 354541 229633 354819
rect 229911 354541 229927 354819
rect 227757 353859 228067 353875
rect 227757 353581 227773 353859
rect 228051 353581 228067 353859
rect 222477 349029 222493 349307
rect 222771 349029 222787 349307
rect 222477 331307 222787 349029
rect 222477 331029 222493 331307
rect 222771 331029 222787 331307
rect 222477 313307 222787 331029
rect 222477 313029 222493 313307
rect 222771 313029 222787 313307
rect 222477 295307 222787 313029
rect 222477 295029 222493 295307
rect 222771 295029 222787 295307
rect 222477 277307 222787 295029
rect 222477 277029 222493 277307
rect 222771 277029 222787 277307
rect 222477 259307 222787 277029
rect 222477 259029 222493 259307
rect 222771 259029 222787 259307
rect 222477 241307 222787 259029
rect 222477 241029 222493 241307
rect 222771 241029 222787 241307
rect 222477 223307 222787 241029
rect 222477 223029 222493 223307
rect 222771 223029 222787 223307
rect 222477 205307 222787 223029
rect 222477 205029 222493 205307
rect 222771 205029 222787 205307
rect 222477 187307 222787 205029
rect 222477 187029 222493 187307
rect 222771 187029 222787 187307
rect 222477 169307 222787 187029
rect 222477 169029 222493 169307
rect 222771 169029 222787 169307
rect 222477 151307 222787 169029
rect 222477 151029 222493 151307
rect 222771 151029 222787 151307
rect 222477 133307 222787 151029
rect 222477 133029 222493 133307
rect 222771 133029 222787 133307
rect 222477 115307 222787 133029
rect 222477 115029 222493 115307
rect 222771 115029 222787 115307
rect 222477 97307 222787 115029
rect 222477 97029 222493 97307
rect 222771 97029 222787 97307
rect 222477 79307 222787 97029
rect 222477 79029 222493 79307
rect 222771 79029 222787 79307
rect 222477 61307 222787 79029
rect 222477 61029 222493 61307
rect 222771 61029 222787 61307
rect 222477 43307 222787 61029
rect 222477 43029 222493 43307
rect 222771 43029 222787 43307
rect 222477 25307 222787 43029
rect 222477 25029 222493 25307
rect 222771 25029 222787 25307
rect 222477 7307 222787 25029
rect 222477 7029 222493 7307
rect 222771 7029 222787 7307
rect 213477 -3811 213493 -3533
rect 213771 -3811 213787 -3533
rect 213477 -3827 213787 -3811
rect 222477 -3053 222787 7029
rect 225897 352899 226207 352915
rect 225897 352621 225913 352899
rect 226191 352621 226207 352899
rect 225897 334727 226207 352621
rect 225897 334449 225913 334727
rect 226191 334449 226207 334727
rect 225897 316727 226207 334449
rect 225897 316449 225913 316727
rect 226191 316449 226207 316727
rect 225897 298727 226207 316449
rect 225897 298449 225913 298727
rect 226191 298449 226207 298727
rect 225897 280727 226207 298449
rect 225897 280449 225913 280727
rect 226191 280449 226207 280727
rect 225897 262727 226207 280449
rect 225897 262449 225913 262727
rect 226191 262449 226207 262727
rect 225897 244727 226207 262449
rect 225897 244449 225913 244727
rect 226191 244449 226207 244727
rect 225897 226727 226207 244449
rect 225897 226449 225913 226727
rect 226191 226449 226207 226727
rect 225897 208727 226207 226449
rect 225897 208449 225913 208727
rect 226191 208449 226207 208727
rect 225897 190727 226207 208449
rect 225897 190449 225913 190727
rect 226191 190449 226207 190727
rect 225897 172727 226207 190449
rect 225897 172449 225913 172727
rect 226191 172449 226207 172727
rect 225897 154727 226207 172449
rect 225897 154449 225913 154727
rect 226191 154449 226207 154727
rect 225897 136727 226207 154449
rect 225897 136449 225913 136727
rect 226191 136449 226207 136727
rect 225897 118727 226207 136449
rect 225897 118449 225913 118727
rect 226191 118449 226207 118727
rect 225897 100727 226207 118449
rect 225897 100449 225913 100727
rect 226191 100449 226207 100727
rect 225897 82727 226207 100449
rect 225897 82449 225913 82727
rect 226191 82449 226207 82727
rect 225897 64727 226207 82449
rect 225897 64449 225913 64727
rect 226191 64449 226207 64727
rect 225897 46727 226207 64449
rect 225897 46449 225913 46727
rect 226191 46449 226207 46727
rect 225897 28727 226207 46449
rect 225897 28449 225913 28727
rect 226191 28449 226207 28727
rect 225897 10727 226207 28449
rect 225897 10449 225913 10727
rect 226191 10449 226207 10727
rect 225897 -653 226207 10449
rect 225897 -931 225913 -653
rect 226191 -931 226207 -653
rect 225897 -947 226207 -931
rect 227757 336587 228067 353581
rect 227757 336309 227773 336587
rect 228051 336309 228067 336587
rect 227757 318587 228067 336309
rect 227757 318309 227773 318587
rect 228051 318309 228067 318587
rect 227757 300587 228067 318309
rect 227757 300309 227773 300587
rect 228051 300309 228067 300587
rect 227757 282587 228067 300309
rect 227757 282309 227773 282587
rect 228051 282309 228067 282587
rect 227757 264587 228067 282309
rect 227757 264309 227773 264587
rect 228051 264309 228067 264587
rect 227757 246587 228067 264309
rect 227757 246309 227773 246587
rect 228051 246309 228067 246587
rect 227757 228587 228067 246309
rect 227757 228309 227773 228587
rect 228051 228309 228067 228587
rect 227757 210587 228067 228309
rect 227757 210309 227773 210587
rect 228051 210309 228067 210587
rect 227757 192587 228067 210309
rect 227757 192309 227773 192587
rect 228051 192309 228067 192587
rect 227757 174587 228067 192309
rect 227757 174309 227773 174587
rect 228051 174309 228067 174587
rect 227757 156587 228067 174309
rect 227757 156309 227773 156587
rect 228051 156309 228067 156587
rect 227757 138587 228067 156309
rect 227757 138309 227773 138587
rect 228051 138309 228067 138587
rect 227757 120587 228067 138309
rect 227757 120309 227773 120587
rect 228051 120309 228067 120587
rect 227757 102587 228067 120309
rect 227757 102309 227773 102587
rect 228051 102309 228067 102587
rect 227757 84587 228067 102309
rect 227757 84309 227773 84587
rect 228051 84309 228067 84587
rect 227757 66587 228067 84309
rect 227757 66309 227773 66587
rect 228051 66309 228067 66587
rect 227757 48587 228067 66309
rect 227757 48309 227773 48587
rect 228051 48309 228067 48587
rect 227757 30587 228067 48309
rect 227757 30309 227773 30587
rect 228051 30309 228067 30587
rect 227757 12587 228067 30309
rect 227757 12309 227773 12587
rect 228051 12309 228067 12587
rect 227757 -1613 228067 12309
rect 227757 -1891 227773 -1613
rect 228051 -1891 228067 -1613
rect 227757 -1907 228067 -1891
rect 229617 338447 229927 354541
rect 229617 338169 229633 338447
rect 229911 338169 229927 338447
rect 229617 320447 229927 338169
rect 229617 320169 229633 320447
rect 229911 320169 229927 320447
rect 229617 302447 229927 320169
rect 229617 302169 229633 302447
rect 229911 302169 229927 302447
rect 229617 284447 229927 302169
rect 229617 284169 229633 284447
rect 229911 284169 229927 284447
rect 229617 266447 229927 284169
rect 229617 266169 229633 266447
rect 229911 266169 229927 266447
rect 229617 248447 229927 266169
rect 229617 248169 229633 248447
rect 229911 248169 229927 248447
rect 229617 230447 229927 248169
rect 229617 230169 229633 230447
rect 229911 230169 229927 230447
rect 229617 212447 229927 230169
rect 229617 212169 229633 212447
rect 229911 212169 229927 212447
rect 229617 194447 229927 212169
rect 229617 194169 229633 194447
rect 229911 194169 229927 194447
rect 229617 176447 229927 194169
rect 229617 176169 229633 176447
rect 229911 176169 229927 176447
rect 229617 158447 229927 176169
rect 229617 158169 229633 158447
rect 229911 158169 229927 158447
rect 229617 140447 229927 158169
rect 229617 140169 229633 140447
rect 229911 140169 229927 140447
rect 229617 122447 229927 140169
rect 229617 122169 229633 122447
rect 229911 122169 229927 122447
rect 229617 104447 229927 122169
rect 229617 104169 229633 104447
rect 229911 104169 229927 104447
rect 229617 86447 229927 104169
rect 229617 86169 229633 86447
rect 229911 86169 229927 86447
rect 229617 68447 229927 86169
rect 229617 68169 229633 68447
rect 229911 68169 229927 68447
rect 229617 50447 229927 68169
rect 229617 50169 229633 50447
rect 229911 50169 229927 50447
rect 229617 32447 229927 50169
rect 229617 32169 229633 32447
rect 229911 32169 229927 32447
rect 229617 14447 229927 32169
rect 229617 14169 229633 14447
rect 229911 14169 229927 14447
rect 229617 -2573 229927 14169
rect 229617 -2851 229633 -2573
rect 229911 -2851 229927 -2573
rect 229617 -2867 229927 -2851
rect 231477 340307 231787 355501
rect 240477 355299 240787 355795
rect 240477 355021 240493 355299
rect 240771 355021 240787 355299
rect 238617 354339 238927 354835
rect 238617 354061 238633 354339
rect 238911 354061 238927 354339
rect 236757 353379 237067 353875
rect 236757 353101 236773 353379
rect 237051 353101 237067 353379
rect 231477 340029 231493 340307
rect 231771 340029 231787 340307
rect 231477 322307 231787 340029
rect 231477 322029 231493 322307
rect 231771 322029 231787 322307
rect 231477 304307 231787 322029
rect 231477 304029 231493 304307
rect 231771 304029 231787 304307
rect 231477 286307 231787 304029
rect 231477 286029 231493 286307
rect 231771 286029 231787 286307
rect 231477 268307 231787 286029
rect 231477 268029 231493 268307
rect 231771 268029 231787 268307
rect 231477 250307 231787 268029
rect 231477 250029 231493 250307
rect 231771 250029 231787 250307
rect 231477 232307 231787 250029
rect 231477 232029 231493 232307
rect 231771 232029 231787 232307
rect 231477 214307 231787 232029
rect 231477 214029 231493 214307
rect 231771 214029 231787 214307
rect 231477 196307 231787 214029
rect 231477 196029 231493 196307
rect 231771 196029 231787 196307
rect 231477 178307 231787 196029
rect 231477 178029 231493 178307
rect 231771 178029 231787 178307
rect 231477 160307 231787 178029
rect 231477 160029 231493 160307
rect 231771 160029 231787 160307
rect 231477 142307 231787 160029
rect 231477 142029 231493 142307
rect 231771 142029 231787 142307
rect 231477 124307 231787 142029
rect 231477 124029 231493 124307
rect 231771 124029 231787 124307
rect 231477 106307 231787 124029
rect 231477 106029 231493 106307
rect 231771 106029 231787 106307
rect 231477 88307 231787 106029
rect 231477 88029 231493 88307
rect 231771 88029 231787 88307
rect 231477 70307 231787 88029
rect 231477 70029 231493 70307
rect 231771 70029 231787 70307
rect 231477 52307 231787 70029
rect 231477 52029 231493 52307
rect 231771 52029 231787 52307
rect 231477 34307 231787 52029
rect 231477 34029 231493 34307
rect 231771 34029 231787 34307
rect 231477 16307 231787 34029
rect 231477 16029 231493 16307
rect 231771 16029 231787 16307
rect 222477 -3331 222493 -3053
rect 222771 -3331 222787 -3053
rect 222477 -3827 222787 -3331
rect 231477 -3533 231787 16029
rect 234897 352419 235207 352915
rect 234897 352141 234913 352419
rect 235191 352141 235207 352419
rect 234897 343727 235207 352141
rect 234897 343449 234913 343727
rect 235191 343449 235207 343727
rect 234897 325727 235207 343449
rect 234897 325449 234913 325727
rect 235191 325449 235207 325727
rect 234897 307727 235207 325449
rect 234897 307449 234913 307727
rect 235191 307449 235207 307727
rect 234897 289727 235207 307449
rect 234897 289449 234913 289727
rect 235191 289449 235207 289727
rect 234897 271727 235207 289449
rect 234897 271449 234913 271727
rect 235191 271449 235207 271727
rect 234897 253727 235207 271449
rect 234897 253449 234913 253727
rect 235191 253449 235207 253727
rect 234897 235727 235207 253449
rect 234897 235449 234913 235727
rect 235191 235449 235207 235727
rect 234897 217727 235207 235449
rect 234897 217449 234913 217727
rect 235191 217449 235207 217727
rect 234897 199727 235207 217449
rect 234897 199449 234913 199727
rect 235191 199449 235207 199727
rect 234897 181727 235207 199449
rect 234897 181449 234913 181727
rect 235191 181449 235207 181727
rect 234897 163727 235207 181449
rect 234897 163449 234913 163727
rect 235191 163449 235207 163727
rect 234897 145727 235207 163449
rect 234897 145449 234913 145727
rect 235191 145449 235207 145727
rect 234897 127727 235207 145449
rect 234897 127449 234913 127727
rect 235191 127449 235207 127727
rect 234897 109727 235207 127449
rect 234897 109449 234913 109727
rect 235191 109449 235207 109727
rect 234897 91727 235207 109449
rect 234897 91449 234913 91727
rect 235191 91449 235207 91727
rect 234897 73727 235207 91449
rect 234897 73449 234913 73727
rect 235191 73449 235207 73727
rect 234897 55727 235207 73449
rect 234897 55449 234913 55727
rect 235191 55449 235207 55727
rect 234897 37727 235207 55449
rect 234897 37449 234913 37727
rect 235191 37449 235207 37727
rect 234897 19727 235207 37449
rect 234897 19449 234913 19727
rect 235191 19449 235207 19727
rect 234897 1727 235207 19449
rect 234897 1449 234913 1727
rect 235191 1449 235207 1727
rect 234897 -173 235207 1449
rect 234897 -451 234913 -173
rect 235191 -451 235207 -173
rect 234897 -947 235207 -451
rect 236757 345587 237067 353101
rect 236757 345309 236773 345587
rect 237051 345309 237067 345587
rect 236757 327587 237067 345309
rect 236757 327309 236773 327587
rect 237051 327309 237067 327587
rect 236757 309587 237067 327309
rect 236757 309309 236773 309587
rect 237051 309309 237067 309587
rect 236757 291587 237067 309309
rect 236757 291309 236773 291587
rect 237051 291309 237067 291587
rect 236757 273587 237067 291309
rect 236757 273309 236773 273587
rect 237051 273309 237067 273587
rect 236757 255587 237067 273309
rect 236757 255309 236773 255587
rect 237051 255309 237067 255587
rect 236757 237587 237067 255309
rect 236757 237309 236773 237587
rect 237051 237309 237067 237587
rect 236757 219587 237067 237309
rect 236757 219309 236773 219587
rect 237051 219309 237067 219587
rect 236757 201587 237067 219309
rect 236757 201309 236773 201587
rect 237051 201309 237067 201587
rect 236757 183587 237067 201309
rect 236757 183309 236773 183587
rect 237051 183309 237067 183587
rect 236757 165587 237067 183309
rect 236757 165309 236773 165587
rect 237051 165309 237067 165587
rect 236757 147587 237067 165309
rect 236757 147309 236773 147587
rect 237051 147309 237067 147587
rect 236757 129587 237067 147309
rect 236757 129309 236773 129587
rect 237051 129309 237067 129587
rect 236757 111587 237067 129309
rect 236757 111309 236773 111587
rect 237051 111309 237067 111587
rect 236757 93587 237067 111309
rect 236757 93309 236773 93587
rect 237051 93309 237067 93587
rect 236757 75587 237067 93309
rect 236757 75309 236773 75587
rect 237051 75309 237067 75587
rect 236757 57587 237067 75309
rect 236757 57309 236773 57587
rect 237051 57309 237067 57587
rect 236757 39587 237067 57309
rect 236757 39309 236773 39587
rect 237051 39309 237067 39587
rect 236757 21587 237067 39309
rect 236757 21309 236773 21587
rect 237051 21309 237067 21587
rect 236757 3587 237067 21309
rect 236757 3309 236773 3587
rect 237051 3309 237067 3587
rect 236757 -1133 237067 3309
rect 236757 -1411 236773 -1133
rect 237051 -1411 237067 -1133
rect 236757 -1907 237067 -1411
rect 238617 347447 238927 354061
rect 238617 347169 238633 347447
rect 238911 347169 238927 347447
rect 238617 329447 238927 347169
rect 238617 329169 238633 329447
rect 238911 329169 238927 329447
rect 238617 311447 238927 329169
rect 238617 311169 238633 311447
rect 238911 311169 238927 311447
rect 238617 293447 238927 311169
rect 238617 293169 238633 293447
rect 238911 293169 238927 293447
rect 238617 275447 238927 293169
rect 238617 275169 238633 275447
rect 238911 275169 238927 275447
rect 238617 257447 238927 275169
rect 238617 257169 238633 257447
rect 238911 257169 238927 257447
rect 238617 239447 238927 257169
rect 238617 239169 238633 239447
rect 238911 239169 238927 239447
rect 238617 221447 238927 239169
rect 238617 221169 238633 221447
rect 238911 221169 238927 221447
rect 238617 203447 238927 221169
rect 238617 203169 238633 203447
rect 238911 203169 238927 203447
rect 238617 185447 238927 203169
rect 238617 185169 238633 185447
rect 238911 185169 238927 185447
rect 238617 167447 238927 185169
rect 238617 167169 238633 167447
rect 238911 167169 238927 167447
rect 238617 149447 238927 167169
rect 238617 149169 238633 149447
rect 238911 149169 238927 149447
rect 238617 131447 238927 149169
rect 238617 131169 238633 131447
rect 238911 131169 238927 131447
rect 238617 113447 238927 131169
rect 238617 113169 238633 113447
rect 238911 113169 238927 113447
rect 238617 95447 238927 113169
rect 238617 95169 238633 95447
rect 238911 95169 238927 95447
rect 238617 77447 238927 95169
rect 238617 77169 238633 77447
rect 238911 77169 238927 77447
rect 238617 59447 238927 77169
rect 238617 59169 238633 59447
rect 238911 59169 238927 59447
rect 238617 41447 238927 59169
rect 238617 41169 238633 41447
rect 238911 41169 238927 41447
rect 238617 23447 238927 41169
rect 238617 23169 238633 23447
rect 238911 23169 238927 23447
rect 238617 5447 238927 23169
rect 238617 5169 238633 5447
rect 238911 5169 238927 5447
rect 238617 -2093 238927 5169
rect 238617 -2371 238633 -2093
rect 238911 -2371 238927 -2093
rect 238617 -2867 238927 -2371
rect 240477 349307 240787 355021
rect 249477 355779 249787 355795
rect 249477 355501 249493 355779
rect 249771 355501 249787 355779
rect 247617 354819 247927 354835
rect 247617 354541 247633 354819
rect 247911 354541 247927 354819
rect 245757 353859 246067 353875
rect 245757 353581 245773 353859
rect 246051 353581 246067 353859
rect 240477 349029 240493 349307
rect 240771 349029 240787 349307
rect 240477 331307 240787 349029
rect 240477 331029 240493 331307
rect 240771 331029 240787 331307
rect 240477 313307 240787 331029
rect 240477 313029 240493 313307
rect 240771 313029 240787 313307
rect 240477 295307 240787 313029
rect 240477 295029 240493 295307
rect 240771 295029 240787 295307
rect 240477 277307 240787 295029
rect 240477 277029 240493 277307
rect 240771 277029 240787 277307
rect 240477 259307 240787 277029
rect 240477 259029 240493 259307
rect 240771 259029 240787 259307
rect 240477 241307 240787 259029
rect 240477 241029 240493 241307
rect 240771 241029 240787 241307
rect 240477 223307 240787 241029
rect 240477 223029 240493 223307
rect 240771 223029 240787 223307
rect 240477 205307 240787 223029
rect 240477 205029 240493 205307
rect 240771 205029 240787 205307
rect 240477 187307 240787 205029
rect 240477 187029 240493 187307
rect 240771 187029 240787 187307
rect 240477 169307 240787 187029
rect 240477 169029 240493 169307
rect 240771 169029 240787 169307
rect 240477 151307 240787 169029
rect 240477 151029 240493 151307
rect 240771 151029 240787 151307
rect 240477 133307 240787 151029
rect 240477 133029 240493 133307
rect 240771 133029 240787 133307
rect 240477 115307 240787 133029
rect 240477 115029 240493 115307
rect 240771 115029 240787 115307
rect 240477 97307 240787 115029
rect 240477 97029 240493 97307
rect 240771 97029 240787 97307
rect 240477 79307 240787 97029
rect 240477 79029 240493 79307
rect 240771 79029 240787 79307
rect 240477 61307 240787 79029
rect 240477 61029 240493 61307
rect 240771 61029 240787 61307
rect 240477 43307 240787 61029
rect 240477 43029 240493 43307
rect 240771 43029 240787 43307
rect 240477 25307 240787 43029
rect 240477 25029 240493 25307
rect 240771 25029 240787 25307
rect 240477 7307 240787 25029
rect 240477 7029 240493 7307
rect 240771 7029 240787 7307
rect 231477 -3811 231493 -3533
rect 231771 -3811 231787 -3533
rect 231477 -3827 231787 -3811
rect 240477 -3053 240787 7029
rect 243897 352899 244207 352915
rect 243897 352621 243913 352899
rect 244191 352621 244207 352899
rect 243897 334727 244207 352621
rect 243897 334449 243913 334727
rect 244191 334449 244207 334727
rect 243897 316727 244207 334449
rect 243897 316449 243913 316727
rect 244191 316449 244207 316727
rect 243897 298727 244207 316449
rect 243897 298449 243913 298727
rect 244191 298449 244207 298727
rect 243897 280727 244207 298449
rect 243897 280449 243913 280727
rect 244191 280449 244207 280727
rect 243897 262727 244207 280449
rect 243897 262449 243913 262727
rect 244191 262449 244207 262727
rect 243897 244727 244207 262449
rect 243897 244449 243913 244727
rect 244191 244449 244207 244727
rect 243897 226727 244207 244449
rect 243897 226449 243913 226727
rect 244191 226449 244207 226727
rect 243897 208727 244207 226449
rect 243897 208449 243913 208727
rect 244191 208449 244207 208727
rect 243897 190727 244207 208449
rect 243897 190449 243913 190727
rect 244191 190449 244207 190727
rect 243897 172727 244207 190449
rect 243897 172449 243913 172727
rect 244191 172449 244207 172727
rect 243897 154727 244207 172449
rect 243897 154449 243913 154727
rect 244191 154449 244207 154727
rect 243897 136727 244207 154449
rect 243897 136449 243913 136727
rect 244191 136449 244207 136727
rect 243897 118727 244207 136449
rect 243897 118449 243913 118727
rect 244191 118449 244207 118727
rect 243897 100727 244207 118449
rect 243897 100449 243913 100727
rect 244191 100449 244207 100727
rect 243897 82727 244207 100449
rect 243897 82449 243913 82727
rect 244191 82449 244207 82727
rect 243897 64727 244207 82449
rect 243897 64449 243913 64727
rect 244191 64449 244207 64727
rect 243897 46727 244207 64449
rect 243897 46449 243913 46727
rect 244191 46449 244207 46727
rect 243897 28727 244207 46449
rect 243897 28449 243913 28727
rect 244191 28449 244207 28727
rect 243897 10727 244207 28449
rect 243897 10449 243913 10727
rect 244191 10449 244207 10727
rect 243897 -653 244207 10449
rect 243897 -931 243913 -653
rect 244191 -931 244207 -653
rect 243897 -947 244207 -931
rect 245757 336587 246067 353581
rect 245757 336309 245773 336587
rect 246051 336309 246067 336587
rect 245757 318587 246067 336309
rect 245757 318309 245773 318587
rect 246051 318309 246067 318587
rect 245757 300587 246067 318309
rect 245757 300309 245773 300587
rect 246051 300309 246067 300587
rect 245757 282587 246067 300309
rect 245757 282309 245773 282587
rect 246051 282309 246067 282587
rect 245757 264587 246067 282309
rect 245757 264309 245773 264587
rect 246051 264309 246067 264587
rect 245757 246587 246067 264309
rect 245757 246309 245773 246587
rect 246051 246309 246067 246587
rect 245757 228587 246067 246309
rect 245757 228309 245773 228587
rect 246051 228309 246067 228587
rect 245757 210587 246067 228309
rect 245757 210309 245773 210587
rect 246051 210309 246067 210587
rect 245757 192587 246067 210309
rect 245757 192309 245773 192587
rect 246051 192309 246067 192587
rect 245757 174587 246067 192309
rect 245757 174309 245773 174587
rect 246051 174309 246067 174587
rect 245757 156587 246067 174309
rect 245757 156309 245773 156587
rect 246051 156309 246067 156587
rect 245757 138587 246067 156309
rect 245757 138309 245773 138587
rect 246051 138309 246067 138587
rect 245757 120587 246067 138309
rect 245757 120309 245773 120587
rect 246051 120309 246067 120587
rect 245757 102587 246067 120309
rect 245757 102309 245773 102587
rect 246051 102309 246067 102587
rect 245757 84587 246067 102309
rect 245757 84309 245773 84587
rect 246051 84309 246067 84587
rect 245757 66587 246067 84309
rect 245757 66309 245773 66587
rect 246051 66309 246067 66587
rect 245757 48587 246067 66309
rect 245757 48309 245773 48587
rect 246051 48309 246067 48587
rect 245757 30587 246067 48309
rect 245757 30309 245773 30587
rect 246051 30309 246067 30587
rect 245757 12587 246067 30309
rect 245757 12309 245773 12587
rect 246051 12309 246067 12587
rect 245757 -1613 246067 12309
rect 245757 -1891 245773 -1613
rect 246051 -1891 246067 -1613
rect 245757 -1907 246067 -1891
rect 247617 338447 247927 354541
rect 247617 338169 247633 338447
rect 247911 338169 247927 338447
rect 247617 320447 247927 338169
rect 247617 320169 247633 320447
rect 247911 320169 247927 320447
rect 247617 302447 247927 320169
rect 247617 302169 247633 302447
rect 247911 302169 247927 302447
rect 247617 284447 247927 302169
rect 247617 284169 247633 284447
rect 247911 284169 247927 284447
rect 247617 266447 247927 284169
rect 247617 266169 247633 266447
rect 247911 266169 247927 266447
rect 247617 248447 247927 266169
rect 247617 248169 247633 248447
rect 247911 248169 247927 248447
rect 247617 230447 247927 248169
rect 247617 230169 247633 230447
rect 247911 230169 247927 230447
rect 247617 212447 247927 230169
rect 247617 212169 247633 212447
rect 247911 212169 247927 212447
rect 247617 194447 247927 212169
rect 247617 194169 247633 194447
rect 247911 194169 247927 194447
rect 247617 176447 247927 194169
rect 247617 176169 247633 176447
rect 247911 176169 247927 176447
rect 247617 158447 247927 176169
rect 247617 158169 247633 158447
rect 247911 158169 247927 158447
rect 247617 140447 247927 158169
rect 247617 140169 247633 140447
rect 247911 140169 247927 140447
rect 247617 122447 247927 140169
rect 247617 122169 247633 122447
rect 247911 122169 247927 122447
rect 247617 104447 247927 122169
rect 247617 104169 247633 104447
rect 247911 104169 247927 104447
rect 247617 86447 247927 104169
rect 247617 86169 247633 86447
rect 247911 86169 247927 86447
rect 247617 68447 247927 86169
rect 247617 68169 247633 68447
rect 247911 68169 247927 68447
rect 247617 50447 247927 68169
rect 247617 50169 247633 50447
rect 247911 50169 247927 50447
rect 247617 32447 247927 50169
rect 247617 32169 247633 32447
rect 247911 32169 247927 32447
rect 247617 14447 247927 32169
rect 247617 14169 247633 14447
rect 247911 14169 247927 14447
rect 247617 -2573 247927 14169
rect 247617 -2851 247633 -2573
rect 247911 -2851 247927 -2573
rect 247617 -2867 247927 -2851
rect 249477 340307 249787 355501
rect 258477 355299 258787 355795
rect 258477 355021 258493 355299
rect 258771 355021 258787 355299
rect 256617 354339 256927 354835
rect 256617 354061 256633 354339
rect 256911 354061 256927 354339
rect 254757 353379 255067 353875
rect 254757 353101 254773 353379
rect 255051 353101 255067 353379
rect 249477 340029 249493 340307
rect 249771 340029 249787 340307
rect 249477 322307 249787 340029
rect 249477 322029 249493 322307
rect 249771 322029 249787 322307
rect 249477 304307 249787 322029
rect 249477 304029 249493 304307
rect 249771 304029 249787 304307
rect 249477 286307 249787 304029
rect 249477 286029 249493 286307
rect 249771 286029 249787 286307
rect 249477 268307 249787 286029
rect 249477 268029 249493 268307
rect 249771 268029 249787 268307
rect 249477 250307 249787 268029
rect 249477 250029 249493 250307
rect 249771 250029 249787 250307
rect 249477 232307 249787 250029
rect 249477 232029 249493 232307
rect 249771 232029 249787 232307
rect 249477 214307 249787 232029
rect 249477 214029 249493 214307
rect 249771 214029 249787 214307
rect 249477 196307 249787 214029
rect 249477 196029 249493 196307
rect 249771 196029 249787 196307
rect 249477 178307 249787 196029
rect 249477 178029 249493 178307
rect 249771 178029 249787 178307
rect 249477 160307 249787 178029
rect 249477 160029 249493 160307
rect 249771 160029 249787 160307
rect 249477 142307 249787 160029
rect 249477 142029 249493 142307
rect 249771 142029 249787 142307
rect 249477 124307 249787 142029
rect 249477 124029 249493 124307
rect 249771 124029 249787 124307
rect 249477 106307 249787 124029
rect 249477 106029 249493 106307
rect 249771 106029 249787 106307
rect 249477 88307 249787 106029
rect 249477 88029 249493 88307
rect 249771 88029 249787 88307
rect 249477 70307 249787 88029
rect 249477 70029 249493 70307
rect 249771 70029 249787 70307
rect 249477 52307 249787 70029
rect 249477 52029 249493 52307
rect 249771 52029 249787 52307
rect 249477 34307 249787 52029
rect 249477 34029 249493 34307
rect 249771 34029 249787 34307
rect 249477 16307 249787 34029
rect 249477 16029 249493 16307
rect 249771 16029 249787 16307
rect 240477 -3331 240493 -3053
rect 240771 -3331 240787 -3053
rect 240477 -3827 240787 -3331
rect 249477 -3533 249787 16029
rect 252897 352419 253207 352915
rect 252897 352141 252913 352419
rect 253191 352141 253207 352419
rect 252897 343727 253207 352141
rect 252897 343449 252913 343727
rect 253191 343449 253207 343727
rect 252897 325727 253207 343449
rect 252897 325449 252913 325727
rect 253191 325449 253207 325727
rect 252897 307727 253207 325449
rect 252897 307449 252913 307727
rect 253191 307449 253207 307727
rect 252897 289727 253207 307449
rect 252897 289449 252913 289727
rect 253191 289449 253207 289727
rect 252897 271727 253207 289449
rect 252897 271449 252913 271727
rect 253191 271449 253207 271727
rect 252897 253727 253207 271449
rect 252897 253449 252913 253727
rect 253191 253449 253207 253727
rect 252897 235727 253207 253449
rect 252897 235449 252913 235727
rect 253191 235449 253207 235727
rect 252897 217727 253207 235449
rect 252897 217449 252913 217727
rect 253191 217449 253207 217727
rect 252897 199727 253207 217449
rect 252897 199449 252913 199727
rect 253191 199449 253207 199727
rect 252897 181727 253207 199449
rect 252897 181449 252913 181727
rect 253191 181449 253207 181727
rect 252897 163727 253207 181449
rect 252897 163449 252913 163727
rect 253191 163449 253207 163727
rect 252897 145727 253207 163449
rect 252897 145449 252913 145727
rect 253191 145449 253207 145727
rect 252897 127727 253207 145449
rect 252897 127449 252913 127727
rect 253191 127449 253207 127727
rect 252897 109727 253207 127449
rect 252897 109449 252913 109727
rect 253191 109449 253207 109727
rect 252897 91727 253207 109449
rect 252897 91449 252913 91727
rect 253191 91449 253207 91727
rect 252897 73727 253207 91449
rect 252897 73449 252913 73727
rect 253191 73449 253207 73727
rect 252897 55727 253207 73449
rect 252897 55449 252913 55727
rect 253191 55449 253207 55727
rect 252897 37727 253207 55449
rect 252897 37449 252913 37727
rect 253191 37449 253207 37727
rect 252897 19727 253207 37449
rect 252897 19449 252913 19727
rect 253191 19449 253207 19727
rect 252897 1727 253207 19449
rect 252897 1449 252913 1727
rect 253191 1449 253207 1727
rect 252897 -173 253207 1449
rect 252897 -451 252913 -173
rect 253191 -451 253207 -173
rect 252897 -947 253207 -451
rect 254757 345587 255067 353101
rect 254757 345309 254773 345587
rect 255051 345309 255067 345587
rect 254757 327587 255067 345309
rect 254757 327309 254773 327587
rect 255051 327309 255067 327587
rect 254757 309587 255067 327309
rect 254757 309309 254773 309587
rect 255051 309309 255067 309587
rect 254757 291587 255067 309309
rect 254757 291309 254773 291587
rect 255051 291309 255067 291587
rect 254757 273587 255067 291309
rect 254757 273309 254773 273587
rect 255051 273309 255067 273587
rect 254757 255587 255067 273309
rect 254757 255309 254773 255587
rect 255051 255309 255067 255587
rect 254757 237587 255067 255309
rect 254757 237309 254773 237587
rect 255051 237309 255067 237587
rect 254757 219587 255067 237309
rect 254757 219309 254773 219587
rect 255051 219309 255067 219587
rect 254757 201587 255067 219309
rect 254757 201309 254773 201587
rect 255051 201309 255067 201587
rect 254757 183587 255067 201309
rect 254757 183309 254773 183587
rect 255051 183309 255067 183587
rect 254757 165587 255067 183309
rect 254757 165309 254773 165587
rect 255051 165309 255067 165587
rect 254757 147587 255067 165309
rect 254757 147309 254773 147587
rect 255051 147309 255067 147587
rect 254757 129587 255067 147309
rect 254757 129309 254773 129587
rect 255051 129309 255067 129587
rect 254757 111587 255067 129309
rect 254757 111309 254773 111587
rect 255051 111309 255067 111587
rect 254757 93587 255067 111309
rect 254757 93309 254773 93587
rect 255051 93309 255067 93587
rect 254757 75587 255067 93309
rect 254757 75309 254773 75587
rect 255051 75309 255067 75587
rect 254757 57587 255067 75309
rect 254757 57309 254773 57587
rect 255051 57309 255067 57587
rect 254757 39587 255067 57309
rect 254757 39309 254773 39587
rect 255051 39309 255067 39587
rect 254757 21587 255067 39309
rect 254757 21309 254773 21587
rect 255051 21309 255067 21587
rect 254757 3587 255067 21309
rect 254757 3309 254773 3587
rect 255051 3309 255067 3587
rect 254757 -1133 255067 3309
rect 254757 -1411 254773 -1133
rect 255051 -1411 255067 -1133
rect 254757 -1907 255067 -1411
rect 256617 347447 256927 354061
rect 256617 347169 256633 347447
rect 256911 347169 256927 347447
rect 256617 329447 256927 347169
rect 256617 329169 256633 329447
rect 256911 329169 256927 329447
rect 256617 311447 256927 329169
rect 256617 311169 256633 311447
rect 256911 311169 256927 311447
rect 256617 293447 256927 311169
rect 256617 293169 256633 293447
rect 256911 293169 256927 293447
rect 256617 275447 256927 293169
rect 256617 275169 256633 275447
rect 256911 275169 256927 275447
rect 256617 257447 256927 275169
rect 256617 257169 256633 257447
rect 256911 257169 256927 257447
rect 256617 239447 256927 257169
rect 256617 239169 256633 239447
rect 256911 239169 256927 239447
rect 256617 221447 256927 239169
rect 256617 221169 256633 221447
rect 256911 221169 256927 221447
rect 256617 203447 256927 221169
rect 256617 203169 256633 203447
rect 256911 203169 256927 203447
rect 256617 185447 256927 203169
rect 256617 185169 256633 185447
rect 256911 185169 256927 185447
rect 256617 167447 256927 185169
rect 256617 167169 256633 167447
rect 256911 167169 256927 167447
rect 256617 149447 256927 167169
rect 256617 149169 256633 149447
rect 256911 149169 256927 149447
rect 256617 131447 256927 149169
rect 256617 131169 256633 131447
rect 256911 131169 256927 131447
rect 256617 113447 256927 131169
rect 256617 113169 256633 113447
rect 256911 113169 256927 113447
rect 256617 95447 256927 113169
rect 256617 95169 256633 95447
rect 256911 95169 256927 95447
rect 256617 77447 256927 95169
rect 256617 77169 256633 77447
rect 256911 77169 256927 77447
rect 256617 59447 256927 77169
rect 256617 59169 256633 59447
rect 256911 59169 256927 59447
rect 256617 41447 256927 59169
rect 256617 41169 256633 41447
rect 256911 41169 256927 41447
rect 256617 23447 256927 41169
rect 256617 23169 256633 23447
rect 256911 23169 256927 23447
rect 256617 5447 256927 23169
rect 256617 5169 256633 5447
rect 256911 5169 256927 5447
rect 256617 -2093 256927 5169
rect 256617 -2371 256633 -2093
rect 256911 -2371 256927 -2093
rect 256617 -2867 256927 -2371
rect 258477 349307 258787 355021
rect 267477 355779 267787 355795
rect 267477 355501 267493 355779
rect 267771 355501 267787 355779
rect 265617 354819 265927 354835
rect 265617 354541 265633 354819
rect 265911 354541 265927 354819
rect 263757 353859 264067 353875
rect 263757 353581 263773 353859
rect 264051 353581 264067 353859
rect 258477 349029 258493 349307
rect 258771 349029 258787 349307
rect 258477 331307 258787 349029
rect 258477 331029 258493 331307
rect 258771 331029 258787 331307
rect 258477 313307 258787 331029
rect 258477 313029 258493 313307
rect 258771 313029 258787 313307
rect 258477 295307 258787 313029
rect 258477 295029 258493 295307
rect 258771 295029 258787 295307
rect 258477 277307 258787 295029
rect 258477 277029 258493 277307
rect 258771 277029 258787 277307
rect 258477 259307 258787 277029
rect 258477 259029 258493 259307
rect 258771 259029 258787 259307
rect 258477 241307 258787 259029
rect 258477 241029 258493 241307
rect 258771 241029 258787 241307
rect 258477 223307 258787 241029
rect 258477 223029 258493 223307
rect 258771 223029 258787 223307
rect 258477 205307 258787 223029
rect 258477 205029 258493 205307
rect 258771 205029 258787 205307
rect 258477 187307 258787 205029
rect 258477 187029 258493 187307
rect 258771 187029 258787 187307
rect 258477 169307 258787 187029
rect 258477 169029 258493 169307
rect 258771 169029 258787 169307
rect 258477 151307 258787 169029
rect 258477 151029 258493 151307
rect 258771 151029 258787 151307
rect 258477 133307 258787 151029
rect 258477 133029 258493 133307
rect 258771 133029 258787 133307
rect 258477 115307 258787 133029
rect 258477 115029 258493 115307
rect 258771 115029 258787 115307
rect 258477 97307 258787 115029
rect 258477 97029 258493 97307
rect 258771 97029 258787 97307
rect 258477 79307 258787 97029
rect 258477 79029 258493 79307
rect 258771 79029 258787 79307
rect 258477 61307 258787 79029
rect 258477 61029 258493 61307
rect 258771 61029 258787 61307
rect 258477 43307 258787 61029
rect 258477 43029 258493 43307
rect 258771 43029 258787 43307
rect 258477 25307 258787 43029
rect 258477 25029 258493 25307
rect 258771 25029 258787 25307
rect 258477 7307 258787 25029
rect 258477 7029 258493 7307
rect 258771 7029 258787 7307
rect 249477 -3811 249493 -3533
rect 249771 -3811 249787 -3533
rect 249477 -3827 249787 -3811
rect 258477 -3053 258787 7029
rect 261897 352899 262207 352915
rect 261897 352621 261913 352899
rect 262191 352621 262207 352899
rect 261897 334727 262207 352621
rect 261897 334449 261913 334727
rect 262191 334449 262207 334727
rect 261897 316727 262207 334449
rect 261897 316449 261913 316727
rect 262191 316449 262207 316727
rect 261897 298727 262207 316449
rect 261897 298449 261913 298727
rect 262191 298449 262207 298727
rect 261897 280727 262207 298449
rect 261897 280449 261913 280727
rect 262191 280449 262207 280727
rect 261897 262727 262207 280449
rect 261897 262449 261913 262727
rect 262191 262449 262207 262727
rect 261897 244727 262207 262449
rect 261897 244449 261913 244727
rect 262191 244449 262207 244727
rect 261897 226727 262207 244449
rect 261897 226449 261913 226727
rect 262191 226449 262207 226727
rect 261897 208727 262207 226449
rect 261897 208449 261913 208727
rect 262191 208449 262207 208727
rect 261897 190727 262207 208449
rect 261897 190449 261913 190727
rect 262191 190449 262207 190727
rect 261897 172727 262207 190449
rect 261897 172449 261913 172727
rect 262191 172449 262207 172727
rect 261897 154727 262207 172449
rect 261897 154449 261913 154727
rect 262191 154449 262207 154727
rect 261897 136727 262207 154449
rect 261897 136449 261913 136727
rect 262191 136449 262207 136727
rect 261897 118727 262207 136449
rect 261897 118449 261913 118727
rect 262191 118449 262207 118727
rect 261897 100727 262207 118449
rect 261897 100449 261913 100727
rect 262191 100449 262207 100727
rect 261897 82727 262207 100449
rect 261897 82449 261913 82727
rect 262191 82449 262207 82727
rect 261897 64727 262207 82449
rect 261897 64449 261913 64727
rect 262191 64449 262207 64727
rect 261897 46727 262207 64449
rect 261897 46449 261913 46727
rect 262191 46449 262207 46727
rect 261897 28727 262207 46449
rect 261897 28449 261913 28727
rect 262191 28449 262207 28727
rect 261897 10727 262207 28449
rect 261897 10449 261913 10727
rect 262191 10449 262207 10727
rect 261897 -653 262207 10449
rect 261897 -931 261913 -653
rect 262191 -931 262207 -653
rect 261897 -947 262207 -931
rect 263757 336587 264067 353581
rect 263757 336309 263773 336587
rect 264051 336309 264067 336587
rect 263757 318587 264067 336309
rect 263757 318309 263773 318587
rect 264051 318309 264067 318587
rect 263757 300587 264067 318309
rect 263757 300309 263773 300587
rect 264051 300309 264067 300587
rect 263757 282587 264067 300309
rect 263757 282309 263773 282587
rect 264051 282309 264067 282587
rect 263757 264587 264067 282309
rect 263757 264309 263773 264587
rect 264051 264309 264067 264587
rect 263757 246587 264067 264309
rect 263757 246309 263773 246587
rect 264051 246309 264067 246587
rect 263757 228587 264067 246309
rect 263757 228309 263773 228587
rect 264051 228309 264067 228587
rect 263757 210587 264067 228309
rect 263757 210309 263773 210587
rect 264051 210309 264067 210587
rect 263757 192587 264067 210309
rect 263757 192309 263773 192587
rect 264051 192309 264067 192587
rect 263757 174587 264067 192309
rect 263757 174309 263773 174587
rect 264051 174309 264067 174587
rect 263757 156587 264067 174309
rect 263757 156309 263773 156587
rect 264051 156309 264067 156587
rect 263757 138587 264067 156309
rect 263757 138309 263773 138587
rect 264051 138309 264067 138587
rect 263757 120587 264067 138309
rect 263757 120309 263773 120587
rect 264051 120309 264067 120587
rect 263757 102587 264067 120309
rect 263757 102309 263773 102587
rect 264051 102309 264067 102587
rect 263757 84587 264067 102309
rect 263757 84309 263773 84587
rect 264051 84309 264067 84587
rect 263757 66587 264067 84309
rect 263757 66309 263773 66587
rect 264051 66309 264067 66587
rect 263757 48587 264067 66309
rect 263757 48309 263773 48587
rect 264051 48309 264067 48587
rect 263757 30587 264067 48309
rect 263757 30309 263773 30587
rect 264051 30309 264067 30587
rect 263757 12587 264067 30309
rect 263757 12309 263773 12587
rect 264051 12309 264067 12587
rect 263757 -1613 264067 12309
rect 263757 -1891 263773 -1613
rect 264051 -1891 264067 -1613
rect 263757 -1907 264067 -1891
rect 265617 338447 265927 354541
rect 265617 338169 265633 338447
rect 265911 338169 265927 338447
rect 265617 320447 265927 338169
rect 265617 320169 265633 320447
rect 265911 320169 265927 320447
rect 265617 302447 265927 320169
rect 265617 302169 265633 302447
rect 265911 302169 265927 302447
rect 265617 284447 265927 302169
rect 265617 284169 265633 284447
rect 265911 284169 265927 284447
rect 265617 266447 265927 284169
rect 265617 266169 265633 266447
rect 265911 266169 265927 266447
rect 265617 248447 265927 266169
rect 265617 248169 265633 248447
rect 265911 248169 265927 248447
rect 265617 230447 265927 248169
rect 265617 230169 265633 230447
rect 265911 230169 265927 230447
rect 265617 212447 265927 230169
rect 265617 212169 265633 212447
rect 265911 212169 265927 212447
rect 265617 194447 265927 212169
rect 265617 194169 265633 194447
rect 265911 194169 265927 194447
rect 265617 176447 265927 194169
rect 265617 176169 265633 176447
rect 265911 176169 265927 176447
rect 265617 158447 265927 176169
rect 265617 158169 265633 158447
rect 265911 158169 265927 158447
rect 265617 140447 265927 158169
rect 265617 140169 265633 140447
rect 265911 140169 265927 140447
rect 265617 122447 265927 140169
rect 265617 122169 265633 122447
rect 265911 122169 265927 122447
rect 265617 104447 265927 122169
rect 265617 104169 265633 104447
rect 265911 104169 265927 104447
rect 265617 86447 265927 104169
rect 265617 86169 265633 86447
rect 265911 86169 265927 86447
rect 265617 68447 265927 86169
rect 265617 68169 265633 68447
rect 265911 68169 265927 68447
rect 265617 50447 265927 68169
rect 265617 50169 265633 50447
rect 265911 50169 265927 50447
rect 265617 32447 265927 50169
rect 265617 32169 265633 32447
rect 265911 32169 265927 32447
rect 265617 14447 265927 32169
rect 265617 14169 265633 14447
rect 265911 14169 265927 14447
rect 265617 -2573 265927 14169
rect 265617 -2851 265633 -2573
rect 265911 -2851 265927 -2573
rect 265617 -2867 265927 -2851
rect 267477 340307 267787 355501
rect 276477 355299 276787 355795
rect 276477 355021 276493 355299
rect 276771 355021 276787 355299
rect 274617 354339 274927 354835
rect 274617 354061 274633 354339
rect 274911 354061 274927 354339
rect 272757 353379 273067 353875
rect 272757 353101 272773 353379
rect 273051 353101 273067 353379
rect 267477 340029 267493 340307
rect 267771 340029 267787 340307
rect 267477 322307 267787 340029
rect 267477 322029 267493 322307
rect 267771 322029 267787 322307
rect 267477 304307 267787 322029
rect 267477 304029 267493 304307
rect 267771 304029 267787 304307
rect 267477 286307 267787 304029
rect 267477 286029 267493 286307
rect 267771 286029 267787 286307
rect 267477 268307 267787 286029
rect 267477 268029 267493 268307
rect 267771 268029 267787 268307
rect 267477 250307 267787 268029
rect 267477 250029 267493 250307
rect 267771 250029 267787 250307
rect 267477 232307 267787 250029
rect 267477 232029 267493 232307
rect 267771 232029 267787 232307
rect 267477 214307 267787 232029
rect 267477 214029 267493 214307
rect 267771 214029 267787 214307
rect 267477 196307 267787 214029
rect 267477 196029 267493 196307
rect 267771 196029 267787 196307
rect 267477 178307 267787 196029
rect 267477 178029 267493 178307
rect 267771 178029 267787 178307
rect 267477 160307 267787 178029
rect 267477 160029 267493 160307
rect 267771 160029 267787 160307
rect 267477 142307 267787 160029
rect 267477 142029 267493 142307
rect 267771 142029 267787 142307
rect 267477 124307 267787 142029
rect 267477 124029 267493 124307
rect 267771 124029 267787 124307
rect 267477 106307 267787 124029
rect 267477 106029 267493 106307
rect 267771 106029 267787 106307
rect 267477 88307 267787 106029
rect 267477 88029 267493 88307
rect 267771 88029 267787 88307
rect 267477 70307 267787 88029
rect 267477 70029 267493 70307
rect 267771 70029 267787 70307
rect 267477 52307 267787 70029
rect 267477 52029 267493 52307
rect 267771 52029 267787 52307
rect 267477 34307 267787 52029
rect 267477 34029 267493 34307
rect 267771 34029 267787 34307
rect 267477 16307 267787 34029
rect 267477 16029 267493 16307
rect 267771 16029 267787 16307
rect 258477 -3331 258493 -3053
rect 258771 -3331 258787 -3053
rect 258477 -3827 258787 -3331
rect 267477 -3533 267787 16029
rect 270897 352419 271207 352915
rect 270897 352141 270913 352419
rect 271191 352141 271207 352419
rect 270897 343727 271207 352141
rect 270897 343449 270913 343727
rect 271191 343449 271207 343727
rect 270897 325727 271207 343449
rect 270897 325449 270913 325727
rect 271191 325449 271207 325727
rect 270897 307727 271207 325449
rect 270897 307449 270913 307727
rect 271191 307449 271207 307727
rect 270897 289727 271207 307449
rect 270897 289449 270913 289727
rect 271191 289449 271207 289727
rect 270897 271727 271207 289449
rect 270897 271449 270913 271727
rect 271191 271449 271207 271727
rect 270897 253727 271207 271449
rect 270897 253449 270913 253727
rect 271191 253449 271207 253727
rect 270897 235727 271207 253449
rect 270897 235449 270913 235727
rect 271191 235449 271207 235727
rect 270897 217727 271207 235449
rect 270897 217449 270913 217727
rect 271191 217449 271207 217727
rect 270897 199727 271207 217449
rect 270897 199449 270913 199727
rect 271191 199449 271207 199727
rect 270897 181727 271207 199449
rect 270897 181449 270913 181727
rect 271191 181449 271207 181727
rect 270897 163727 271207 181449
rect 270897 163449 270913 163727
rect 271191 163449 271207 163727
rect 270897 145727 271207 163449
rect 270897 145449 270913 145727
rect 271191 145449 271207 145727
rect 270897 127727 271207 145449
rect 270897 127449 270913 127727
rect 271191 127449 271207 127727
rect 270897 109727 271207 127449
rect 270897 109449 270913 109727
rect 271191 109449 271207 109727
rect 270897 91727 271207 109449
rect 270897 91449 270913 91727
rect 271191 91449 271207 91727
rect 270897 73727 271207 91449
rect 270897 73449 270913 73727
rect 271191 73449 271207 73727
rect 270897 55727 271207 73449
rect 270897 55449 270913 55727
rect 271191 55449 271207 55727
rect 270897 37727 271207 55449
rect 270897 37449 270913 37727
rect 271191 37449 271207 37727
rect 270897 19727 271207 37449
rect 270897 19449 270913 19727
rect 271191 19449 271207 19727
rect 270897 1727 271207 19449
rect 270897 1449 270913 1727
rect 271191 1449 271207 1727
rect 270897 -173 271207 1449
rect 270897 -451 270913 -173
rect 271191 -451 271207 -173
rect 270897 -947 271207 -451
rect 272757 345587 273067 353101
rect 272757 345309 272773 345587
rect 273051 345309 273067 345587
rect 272757 327587 273067 345309
rect 272757 327309 272773 327587
rect 273051 327309 273067 327587
rect 272757 309587 273067 327309
rect 272757 309309 272773 309587
rect 273051 309309 273067 309587
rect 272757 291587 273067 309309
rect 272757 291309 272773 291587
rect 273051 291309 273067 291587
rect 272757 273587 273067 291309
rect 272757 273309 272773 273587
rect 273051 273309 273067 273587
rect 272757 255587 273067 273309
rect 272757 255309 272773 255587
rect 273051 255309 273067 255587
rect 272757 237587 273067 255309
rect 272757 237309 272773 237587
rect 273051 237309 273067 237587
rect 272757 219587 273067 237309
rect 272757 219309 272773 219587
rect 273051 219309 273067 219587
rect 272757 201587 273067 219309
rect 272757 201309 272773 201587
rect 273051 201309 273067 201587
rect 272757 183587 273067 201309
rect 272757 183309 272773 183587
rect 273051 183309 273067 183587
rect 272757 165587 273067 183309
rect 272757 165309 272773 165587
rect 273051 165309 273067 165587
rect 272757 147587 273067 165309
rect 272757 147309 272773 147587
rect 273051 147309 273067 147587
rect 272757 129587 273067 147309
rect 272757 129309 272773 129587
rect 273051 129309 273067 129587
rect 272757 111587 273067 129309
rect 272757 111309 272773 111587
rect 273051 111309 273067 111587
rect 272757 93587 273067 111309
rect 272757 93309 272773 93587
rect 273051 93309 273067 93587
rect 272757 75587 273067 93309
rect 272757 75309 272773 75587
rect 273051 75309 273067 75587
rect 272757 57587 273067 75309
rect 272757 57309 272773 57587
rect 273051 57309 273067 57587
rect 272757 39587 273067 57309
rect 272757 39309 272773 39587
rect 273051 39309 273067 39587
rect 272757 21587 273067 39309
rect 272757 21309 272773 21587
rect 273051 21309 273067 21587
rect 272757 3587 273067 21309
rect 272757 3309 272773 3587
rect 273051 3309 273067 3587
rect 272757 -1133 273067 3309
rect 272757 -1411 272773 -1133
rect 273051 -1411 273067 -1133
rect 272757 -1907 273067 -1411
rect 274617 347447 274927 354061
rect 274617 347169 274633 347447
rect 274911 347169 274927 347447
rect 274617 329447 274927 347169
rect 274617 329169 274633 329447
rect 274911 329169 274927 329447
rect 274617 311447 274927 329169
rect 274617 311169 274633 311447
rect 274911 311169 274927 311447
rect 274617 293447 274927 311169
rect 274617 293169 274633 293447
rect 274911 293169 274927 293447
rect 274617 275447 274927 293169
rect 274617 275169 274633 275447
rect 274911 275169 274927 275447
rect 274617 257447 274927 275169
rect 274617 257169 274633 257447
rect 274911 257169 274927 257447
rect 274617 239447 274927 257169
rect 274617 239169 274633 239447
rect 274911 239169 274927 239447
rect 274617 221447 274927 239169
rect 274617 221169 274633 221447
rect 274911 221169 274927 221447
rect 274617 203447 274927 221169
rect 274617 203169 274633 203447
rect 274911 203169 274927 203447
rect 274617 185447 274927 203169
rect 274617 185169 274633 185447
rect 274911 185169 274927 185447
rect 274617 167447 274927 185169
rect 274617 167169 274633 167447
rect 274911 167169 274927 167447
rect 274617 149447 274927 167169
rect 274617 149169 274633 149447
rect 274911 149169 274927 149447
rect 274617 131447 274927 149169
rect 274617 131169 274633 131447
rect 274911 131169 274927 131447
rect 274617 113447 274927 131169
rect 274617 113169 274633 113447
rect 274911 113169 274927 113447
rect 274617 95447 274927 113169
rect 274617 95169 274633 95447
rect 274911 95169 274927 95447
rect 274617 77447 274927 95169
rect 274617 77169 274633 77447
rect 274911 77169 274927 77447
rect 274617 59447 274927 77169
rect 274617 59169 274633 59447
rect 274911 59169 274927 59447
rect 274617 41447 274927 59169
rect 274617 41169 274633 41447
rect 274911 41169 274927 41447
rect 274617 23447 274927 41169
rect 274617 23169 274633 23447
rect 274911 23169 274927 23447
rect 274617 5447 274927 23169
rect 274617 5169 274633 5447
rect 274911 5169 274927 5447
rect 274617 -2093 274927 5169
rect 274617 -2371 274633 -2093
rect 274911 -2371 274927 -2093
rect 274617 -2867 274927 -2371
rect 276477 349307 276787 355021
rect 285477 355779 285787 355795
rect 285477 355501 285493 355779
rect 285771 355501 285787 355779
rect 283617 354819 283927 354835
rect 283617 354541 283633 354819
rect 283911 354541 283927 354819
rect 281757 353859 282067 353875
rect 281757 353581 281773 353859
rect 282051 353581 282067 353859
rect 276477 349029 276493 349307
rect 276771 349029 276787 349307
rect 276477 331307 276787 349029
rect 276477 331029 276493 331307
rect 276771 331029 276787 331307
rect 276477 313307 276787 331029
rect 276477 313029 276493 313307
rect 276771 313029 276787 313307
rect 276477 295307 276787 313029
rect 276477 295029 276493 295307
rect 276771 295029 276787 295307
rect 276477 277307 276787 295029
rect 276477 277029 276493 277307
rect 276771 277029 276787 277307
rect 276477 259307 276787 277029
rect 276477 259029 276493 259307
rect 276771 259029 276787 259307
rect 276477 241307 276787 259029
rect 276477 241029 276493 241307
rect 276771 241029 276787 241307
rect 276477 223307 276787 241029
rect 276477 223029 276493 223307
rect 276771 223029 276787 223307
rect 276477 205307 276787 223029
rect 276477 205029 276493 205307
rect 276771 205029 276787 205307
rect 276477 187307 276787 205029
rect 276477 187029 276493 187307
rect 276771 187029 276787 187307
rect 276477 169307 276787 187029
rect 276477 169029 276493 169307
rect 276771 169029 276787 169307
rect 276477 151307 276787 169029
rect 276477 151029 276493 151307
rect 276771 151029 276787 151307
rect 276477 133307 276787 151029
rect 276477 133029 276493 133307
rect 276771 133029 276787 133307
rect 276477 115307 276787 133029
rect 276477 115029 276493 115307
rect 276771 115029 276787 115307
rect 276477 97307 276787 115029
rect 276477 97029 276493 97307
rect 276771 97029 276787 97307
rect 276477 79307 276787 97029
rect 276477 79029 276493 79307
rect 276771 79029 276787 79307
rect 276477 61307 276787 79029
rect 276477 61029 276493 61307
rect 276771 61029 276787 61307
rect 276477 43307 276787 61029
rect 276477 43029 276493 43307
rect 276771 43029 276787 43307
rect 276477 25307 276787 43029
rect 276477 25029 276493 25307
rect 276771 25029 276787 25307
rect 276477 7307 276787 25029
rect 276477 7029 276493 7307
rect 276771 7029 276787 7307
rect 267477 -3811 267493 -3533
rect 267771 -3811 267787 -3533
rect 267477 -3827 267787 -3811
rect 276477 -3053 276787 7029
rect 279897 352899 280207 352915
rect 279897 352621 279913 352899
rect 280191 352621 280207 352899
rect 279897 334727 280207 352621
rect 279897 334449 279913 334727
rect 280191 334449 280207 334727
rect 279897 316727 280207 334449
rect 279897 316449 279913 316727
rect 280191 316449 280207 316727
rect 279897 298727 280207 316449
rect 279897 298449 279913 298727
rect 280191 298449 280207 298727
rect 279897 280727 280207 298449
rect 279897 280449 279913 280727
rect 280191 280449 280207 280727
rect 279897 262727 280207 280449
rect 279897 262449 279913 262727
rect 280191 262449 280207 262727
rect 279897 244727 280207 262449
rect 279897 244449 279913 244727
rect 280191 244449 280207 244727
rect 279897 226727 280207 244449
rect 279897 226449 279913 226727
rect 280191 226449 280207 226727
rect 279897 208727 280207 226449
rect 279897 208449 279913 208727
rect 280191 208449 280207 208727
rect 279897 190727 280207 208449
rect 279897 190449 279913 190727
rect 280191 190449 280207 190727
rect 279897 172727 280207 190449
rect 279897 172449 279913 172727
rect 280191 172449 280207 172727
rect 279897 154727 280207 172449
rect 279897 154449 279913 154727
rect 280191 154449 280207 154727
rect 279897 136727 280207 154449
rect 279897 136449 279913 136727
rect 280191 136449 280207 136727
rect 279897 118727 280207 136449
rect 279897 118449 279913 118727
rect 280191 118449 280207 118727
rect 279897 100727 280207 118449
rect 279897 100449 279913 100727
rect 280191 100449 280207 100727
rect 279897 82727 280207 100449
rect 279897 82449 279913 82727
rect 280191 82449 280207 82727
rect 279897 64727 280207 82449
rect 279897 64449 279913 64727
rect 280191 64449 280207 64727
rect 279897 46727 280207 64449
rect 279897 46449 279913 46727
rect 280191 46449 280207 46727
rect 279897 28727 280207 46449
rect 279897 28449 279913 28727
rect 280191 28449 280207 28727
rect 279897 10727 280207 28449
rect 279897 10449 279913 10727
rect 280191 10449 280207 10727
rect 279897 -653 280207 10449
rect 279897 -931 279913 -653
rect 280191 -931 280207 -653
rect 279897 -947 280207 -931
rect 281757 336587 282067 353581
rect 281757 336309 281773 336587
rect 282051 336309 282067 336587
rect 281757 318587 282067 336309
rect 281757 318309 281773 318587
rect 282051 318309 282067 318587
rect 281757 300587 282067 318309
rect 281757 300309 281773 300587
rect 282051 300309 282067 300587
rect 281757 282587 282067 300309
rect 281757 282309 281773 282587
rect 282051 282309 282067 282587
rect 281757 264587 282067 282309
rect 281757 264309 281773 264587
rect 282051 264309 282067 264587
rect 281757 246587 282067 264309
rect 281757 246309 281773 246587
rect 282051 246309 282067 246587
rect 281757 228587 282067 246309
rect 281757 228309 281773 228587
rect 282051 228309 282067 228587
rect 281757 210587 282067 228309
rect 281757 210309 281773 210587
rect 282051 210309 282067 210587
rect 281757 192587 282067 210309
rect 281757 192309 281773 192587
rect 282051 192309 282067 192587
rect 281757 174587 282067 192309
rect 281757 174309 281773 174587
rect 282051 174309 282067 174587
rect 281757 156587 282067 174309
rect 281757 156309 281773 156587
rect 282051 156309 282067 156587
rect 281757 138587 282067 156309
rect 281757 138309 281773 138587
rect 282051 138309 282067 138587
rect 281757 120587 282067 138309
rect 281757 120309 281773 120587
rect 282051 120309 282067 120587
rect 281757 102587 282067 120309
rect 281757 102309 281773 102587
rect 282051 102309 282067 102587
rect 281757 84587 282067 102309
rect 281757 84309 281773 84587
rect 282051 84309 282067 84587
rect 281757 66587 282067 84309
rect 281757 66309 281773 66587
rect 282051 66309 282067 66587
rect 281757 48587 282067 66309
rect 281757 48309 281773 48587
rect 282051 48309 282067 48587
rect 281757 30587 282067 48309
rect 281757 30309 281773 30587
rect 282051 30309 282067 30587
rect 281757 12587 282067 30309
rect 281757 12309 281773 12587
rect 282051 12309 282067 12587
rect 281757 -1613 282067 12309
rect 281757 -1891 281773 -1613
rect 282051 -1891 282067 -1613
rect 281757 -1907 282067 -1891
rect 283617 338447 283927 354541
rect 283617 338169 283633 338447
rect 283911 338169 283927 338447
rect 283617 320447 283927 338169
rect 283617 320169 283633 320447
rect 283911 320169 283927 320447
rect 283617 302447 283927 320169
rect 283617 302169 283633 302447
rect 283911 302169 283927 302447
rect 283617 284447 283927 302169
rect 283617 284169 283633 284447
rect 283911 284169 283927 284447
rect 283617 266447 283927 284169
rect 283617 266169 283633 266447
rect 283911 266169 283927 266447
rect 283617 248447 283927 266169
rect 283617 248169 283633 248447
rect 283911 248169 283927 248447
rect 283617 230447 283927 248169
rect 283617 230169 283633 230447
rect 283911 230169 283927 230447
rect 283617 212447 283927 230169
rect 283617 212169 283633 212447
rect 283911 212169 283927 212447
rect 283617 194447 283927 212169
rect 283617 194169 283633 194447
rect 283911 194169 283927 194447
rect 283617 176447 283927 194169
rect 283617 176169 283633 176447
rect 283911 176169 283927 176447
rect 283617 158447 283927 176169
rect 283617 158169 283633 158447
rect 283911 158169 283927 158447
rect 283617 140447 283927 158169
rect 283617 140169 283633 140447
rect 283911 140169 283927 140447
rect 283617 122447 283927 140169
rect 283617 122169 283633 122447
rect 283911 122169 283927 122447
rect 283617 104447 283927 122169
rect 283617 104169 283633 104447
rect 283911 104169 283927 104447
rect 283617 86447 283927 104169
rect 283617 86169 283633 86447
rect 283911 86169 283927 86447
rect 283617 68447 283927 86169
rect 283617 68169 283633 68447
rect 283911 68169 283927 68447
rect 283617 50447 283927 68169
rect 283617 50169 283633 50447
rect 283911 50169 283927 50447
rect 283617 32447 283927 50169
rect 283617 32169 283633 32447
rect 283911 32169 283927 32447
rect 283617 14447 283927 32169
rect 283617 14169 283633 14447
rect 283911 14169 283927 14447
rect 283617 -2573 283927 14169
rect 283617 -2851 283633 -2573
rect 283911 -2851 283927 -2573
rect 283617 -2867 283927 -2851
rect 285477 340307 285787 355501
rect 296015 355779 296325 355795
rect 296015 355501 296031 355779
rect 296309 355501 296325 355779
rect 295535 355299 295845 355315
rect 295535 355021 295551 355299
rect 295829 355021 295845 355299
rect 295055 354819 295365 354835
rect 295055 354541 295071 354819
rect 295349 354541 295365 354819
rect 294575 354339 294885 354355
rect 294575 354061 294591 354339
rect 294869 354061 294885 354339
rect 290757 353379 291067 353875
rect 294095 353859 294405 353875
rect 294095 353581 294111 353859
rect 294389 353581 294405 353859
rect 290757 353101 290773 353379
rect 291051 353101 291067 353379
rect 285477 340029 285493 340307
rect 285771 340029 285787 340307
rect 285477 322307 285787 340029
rect 285477 322029 285493 322307
rect 285771 322029 285787 322307
rect 285477 304307 285787 322029
rect 285477 304029 285493 304307
rect 285771 304029 285787 304307
rect 285477 286307 285787 304029
rect 285477 286029 285493 286307
rect 285771 286029 285787 286307
rect 285477 268307 285787 286029
rect 285477 268029 285493 268307
rect 285771 268029 285787 268307
rect 285477 250307 285787 268029
rect 285477 250029 285493 250307
rect 285771 250029 285787 250307
rect 285477 232307 285787 250029
rect 285477 232029 285493 232307
rect 285771 232029 285787 232307
rect 285477 214307 285787 232029
rect 285477 214029 285493 214307
rect 285771 214029 285787 214307
rect 285477 196307 285787 214029
rect 285477 196029 285493 196307
rect 285771 196029 285787 196307
rect 285477 178307 285787 196029
rect 285477 178029 285493 178307
rect 285771 178029 285787 178307
rect 285477 160307 285787 178029
rect 285477 160029 285493 160307
rect 285771 160029 285787 160307
rect 285477 142307 285787 160029
rect 285477 142029 285493 142307
rect 285771 142029 285787 142307
rect 285477 124307 285787 142029
rect 285477 124029 285493 124307
rect 285771 124029 285787 124307
rect 285477 106307 285787 124029
rect 285477 106029 285493 106307
rect 285771 106029 285787 106307
rect 285477 88307 285787 106029
rect 285477 88029 285493 88307
rect 285771 88029 285787 88307
rect 285477 70307 285787 88029
rect 285477 70029 285493 70307
rect 285771 70029 285787 70307
rect 285477 52307 285787 70029
rect 285477 52029 285493 52307
rect 285771 52029 285787 52307
rect 285477 34307 285787 52029
rect 285477 34029 285493 34307
rect 285771 34029 285787 34307
rect 285477 16307 285787 34029
rect 285477 16029 285493 16307
rect 285771 16029 285787 16307
rect 276477 -3331 276493 -3053
rect 276771 -3331 276787 -3053
rect 276477 -3827 276787 -3331
rect 285477 -3533 285787 16029
rect 288897 352419 289207 352915
rect 288897 352141 288913 352419
rect 289191 352141 289207 352419
rect 288897 343727 289207 352141
rect 288897 343449 288913 343727
rect 289191 343449 289207 343727
rect 288897 325727 289207 343449
rect 288897 325449 288913 325727
rect 289191 325449 289207 325727
rect 288897 307727 289207 325449
rect 288897 307449 288913 307727
rect 289191 307449 289207 307727
rect 288897 289727 289207 307449
rect 288897 289449 288913 289727
rect 289191 289449 289207 289727
rect 288897 271727 289207 289449
rect 288897 271449 288913 271727
rect 289191 271449 289207 271727
rect 288897 253727 289207 271449
rect 288897 253449 288913 253727
rect 289191 253449 289207 253727
rect 288897 235727 289207 253449
rect 288897 235449 288913 235727
rect 289191 235449 289207 235727
rect 288897 217727 289207 235449
rect 288897 217449 288913 217727
rect 289191 217449 289207 217727
rect 288897 199727 289207 217449
rect 288897 199449 288913 199727
rect 289191 199449 289207 199727
rect 288897 181727 289207 199449
rect 288897 181449 288913 181727
rect 289191 181449 289207 181727
rect 288897 163727 289207 181449
rect 288897 163449 288913 163727
rect 289191 163449 289207 163727
rect 288897 145727 289207 163449
rect 288897 145449 288913 145727
rect 289191 145449 289207 145727
rect 288897 127727 289207 145449
rect 288897 127449 288913 127727
rect 289191 127449 289207 127727
rect 288897 109727 289207 127449
rect 288897 109449 288913 109727
rect 289191 109449 289207 109727
rect 288897 91727 289207 109449
rect 288897 91449 288913 91727
rect 289191 91449 289207 91727
rect 288897 73727 289207 91449
rect 288897 73449 288913 73727
rect 289191 73449 289207 73727
rect 288897 55727 289207 73449
rect 288897 55449 288913 55727
rect 289191 55449 289207 55727
rect 288897 37727 289207 55449
rect 288897 37449 288913 37727
rect 289191 37449 289207 37727
rect 288897 19727 289207 37449
rect 288897 19449 288913 19727
rect 289191 19449 289207 19727
rect 288897 1727 289207 19449
rect 288897 1449 288913 1727
rect 289191 1449 289207 1727
rect 288897 -173 289207 1449
rect 288897 -451 288913 -173
rect 289191 -451 289207 -173
rect 288897 -947 289207 -451
rect 290757 345587 291067 353101
rect 293615 353379 293925 353395
rect 293615 353101 293631 353379
rect 293909 353101 293925 353379
rect 293135 352899 293445 352915
rect 293135 352621 293151 352899
rect 293429 352621 293445 352899
rect 290757 345309 290773 345587
rect 291051 345309 291067 345587
rect 290757 327587 291067 345309
rect 290757 327309 290773 327587
rect 291051 327309 291067 327587
rect 290757 309587 291067 327309
rect 290757 309309 290773 309587
rect 291051 309309 291067 309587
rect 290757 291587 291067 309309
rect 290757 291309 290773 291587
rect 291051 291309 291067 291587
rect 290757 273587 291067 291309
rect 290757 273309 290773 273587
rect 291051 273309 291067 273587
rect 290757 255587 291067 273309
rect 290757 255309 290773 255587
rect 291051 255309 291067 255587
rect 290757 237587 291067 255309
rect 290757 237309 290773 237587
rect 291051 237309 291067 237587
rect 290757 219587 291067 237309
rect 290757 219309 290773 219587
rect 291051 219309 291067 219587
rect 290757 201587 291067 219309
rect 290757 201309 290773 201587
rect 291051 201309 291067 201587
rect 290757 183587 291067 201309
rect 290757 183309 290773 183587
rect 291051 183309 291067 183587
rect 290757 165587 291067 183309
rect 290757 165309 290773 165587
rect 291051 165309 291067 165587
rect 290757 147587 291067 165309
rect 290757 147309 290773 147587
rect 291051 147309 291067 147587
rect 290757 129587 291067 147309
rect 290757 129309 290773 129587
rect 291051 129309 291067 129587
rect 290757 111587 291067 129309
rect 290757 111309 290773 111587
rect 291051 111309 291067 111587
rect 290757 93587 291067 111309
rect 290757 93309 290773 93587
rect 291051 93309 291067 93587
rect 290757 75587 291067 93309
rect 290757 75309 290773 75587
rect 291051 75309 291067 75587
rect 290757 57587 291067 75309
rect 290757 57309 290773 57587
rect 291051 57309 291067 57587
rect 290757 39587 291067 57309
rect 290757 39309 290773 39587
rect 291051 39309 291067 39587
rect 290757 21587 291067 39309
rect 290757 21309 290773 21587
rect 291051 21309 291067 21587
rect 290757 3587 291067 21309
rect 290757 3309 290773 3587
rect 291051 3309 291067 3587
rect 290757 -1133 291067 3309
rect 292655 352419 292965 352435
rect 292655 352141 292671 352419
rect 292949 352141 292965 352419
rect 292655 343727 292965 352141
rect 292655 343449 292671 343727
rect 292949 343449 292965 343727
rect 292655 325727 292965 343449
rect 292655 325449 292671 325727
rect 292949 325449 292965 325727
rect 292655 307727 292965 325449
rect 292655 307449 292671 307727
rect 292949 307449 292965 307727
rect 292655 289727 292965 307449
rect 292655 289449 292671 289727
rect 292949 289449 292965 289727
rect 292655 271727 292965 289449
rect 292655 271449 292671 271727
rect 292949 271449 292965 271727
rect 292655 253727 292965 271449
rect 292655 253449 292671 253727
rect 292949 253449 292965 253727
rect 292655 235727 292965 253449
rect 292655 235449 292671 235727
rect 292949 235449 292965 235727
rect 292655 217727 292965 235449
rect 292655 217449 292671 217727
rect 292949 217449 292965 217727
rect 292655 199727 292965 217449
rect 292655 199449 292671 199727
rect 292949 199449 292965 199727
rect 292655 181727 292965 199449
rect 292655 181449 292671 181727
rect 292949 181449 292965 181727
rect 292655 163727 292965 181449
rect 292655 163449 292671 163727
rect 292949 163449 292965 163727
rect 292655 145727 292965 163449
rect 292655 145449 292671 145727
rect 292949 145449 292965 145727
rect 292655 127727 292965 145449
rect 292655 127449 292671 127727
rect 292949 127449 292965 127727
rect 292655 109727 292965 127449
rect 292655 109449 292671 109727
rect 292949 109449 292965 109727
rect 292655 91727 292965 109449
rect 292655 91449 292671 91727
rect 292949 91449 292965 91727
rect 292655 73727 292965 91449
rect 292655 73449 292671 73727
rect 292949 73449 292965 73727
rect 292655 55727 292965 73449
rect 292655 55449 292671 55727
rect 292949 55449 292965 55727
rect 292655 37727 292965 55449
rect 292655 37449 292671 37727
rect 292949 37449 292965 37727
rect 292655 19727 292965 37449
rect 292655 19449 292671 19727
rect 292949 19449 292965 19727
rect 292655 1727 292965 19449
rect 292655 1449 292671 1727
rect 292949 1449 292965 1727
rect 292655 -173 292965 1449
rect 292655 -451 292671 -173
rect 292949 -451 292965 -173
rect 292655 -467 292965 -451
rect 293135 334727 293445 352621
rect 293135 334449 293151 334727
rect 293429 334449 293445 334727
rect 293135 316727 293445 334449
rect 293135 316449 293151 316727
rect 293429 316449 293445 316727
rect 293135 298727 293445 316449
rect 293135 298449 293151 298727
rect 293429 298449 293445 298727
rect 293135 280727 293445 298449
rect 293135 280449 293151 280727
rect 293429 280449 293445 280727
rect 293135 262727 293445 280449
rect 293135 262449 293151 262727
rect 293429 262449 293445 262727
rect 293135 244727 293445 262449
rect 293135 244449 293151 244727
rect 293429 244449 293445 244727
rect 293135 226727 293445 244449
rect 293135 226449 293151 226727
rect 293429 226449 293445 226727
rect 293135 208727 293445 226449
rect 293135 208449 293151 208727
rect 293429 208449 293445 208727
rect 293135 190727 293445 208449
rect 293135 190449 293151 190727
rect 293429 190449 293445 190727
rect 293135 172727 293445 190449
rect 293135 172449 293151 172727
rect 293429 172449 293445 172727
rect 293135 154727 293445 172449
rect 293135 154449 293151 154727
rect 293429 154449 293445 154727
rect 293135 136727 293445 154449
rect 293135 136449 293151 136727
rect 293429 136449 293445 136727
rect 293135 118727 293445 136449
rect 293135 118449 293151 118727
rect 293429 118449 293445 118727
rect 293135 100727 293445 118449
rect 293135 100449 293151 100727
rect 293429 100449 293445 100727
rect 293135 82727 293445 100449
rect 293135 82449 293151 82727
rect 293429 82449 293445 82727
rect 293135 64727 293445 82449
rect 293135 64449 293151 64727
rect 293429 64449 293445 64727
rect 293135 46727 293445 64449
rect 293135 46449 293151 46727
rect 293429 46449 293445 46727
rect 293135 28727 293445 46449
rect 293135 28449 293151 28727
rect 293429 28449 293445 28727
rect 293135 10727 293445 28449
rect 293135 10449 293151 10727
rect 293429 10449 293445 10727
rect 293135 -653 293445 10449
rect 293135 -931 293151 -653
rect 293429 -931 293445 -653
rect 293135 -947 293445 -931
rect 293615 345587 293925 353101
rect 293615 345309 293631 345587
rect 293909 345309 293925 345587
rect 293615 327587 293925 345309
rect 293615 327309 293631 327587
rect 293909 327309 293925 327587
rect 293615 309587 293925 327309
rect 293615 309309 293631 309587
rect 293909 309309 293925 309587
rect 293615 291587 293925 309309
rect 293615 291309 293631 291587
rect 293909 291309 293925 291587
rect 293615 273587 293925 291309
rect 293615 273309 293631 273587
rect 293909 273309 293925 273587
rect 293615 255587 293925 273309
rect 293615 255309 293631 255587
rect 293909 255309 293925 255587
rect 293615 237587 293925 255309
rect 293615 237309 293631 237587
rect 293909 237309 293925 237587
rect 293615 219587 293925 237309
rect 293615 219309 293631 219587
rect 293909 219309 293925 219587
rect 293615 201587 293925 219309
rect 293615 201309 293631 201587
rect 293909 201309 293925 201587
rect 293615 183587 293925 201309
rect 293615 183309 293631 183587
rect 293909 183309 293925 183587
rect 293615 165587 293925 183309
rect 293615 165309 293631 165587
rect 293909 165309 293925 165587
rect 293615 147587 293925 165309
rect 293615 147309 293631 147587
rect 293909 147309 293925 147587
rect 293615 129587 293925 147309
rect 293615 129309 293631 129587
rect 293909 129309 293925 129587
rect 293615 111587 293925 129309
rect 293615 111309 293631 111587
rect 293909 111309 293925 111587
rect 293615 93587 293925 111309
rect 293615 93309 293631 93587
rect 293909 93309 293925 93587
rect 293615 75587 293925 93309
rect 293615 75309 293631 75587
rect 293909 75309 293925 75587
rect 293615 57587 293925 75309
rect 293615 57309 293631 57587
rect 293909 57309 293925 57587
rect 293615 39587 293925 57309
rect 293615 39309 293631 39587
rect 293909 39309 293925 39587
rect 293615 21587 293925 39309
rect 293615 21309 293631 21587
rect 293909 21309 293925 21587
rect 293615 3587 293925 21309
rect 293615 3309 293631 3587
rect 293909 3309 293925 3587
rect 290757 -1411 290773 -1133
rect 291051 -1411 291067 -1133
rect 290757 -1907 291067 -1411
rect 293615 -1133 293925 3309
rect 293615 -1411 293631 -1133
rect 293909 -1411 293925 -1133
rect 293615 -1427 293925 -1411
rect 294095 336587 294405 353581
rect 294095 336309 294111 336587
rect 294389 336309 294405 336587
rect 294095 318587 294405 336309
rect 294095 318309 294111 318587
rect 294389 318309 294405 318587
rect 294095 300587 294405 318309
rect 294095 300309 294111 300587
rect 294389 300309 294405 300587
rect 294095 282587 294405 300309
rect 294095 282309 294111 282587
rect 294389 282309 294405 282587
rect 294095 264587 294405 282309
rect 294095 264309 294111 264587
rect 294389 264309 294405 264587
rect 294095 246587 294405 264309
rect 294095 246309 294111 246587
rect 294389 246309 294405 246587
rect 294095 228587 294405 246309
rect 294095 228309 294111 228587
rect 294389 228309 294405 228587
rect 294095 210587 294405 228309
rect 294095 210309 294111 210587
rect 294389 210309 294405 210587
rect 294095 192587 294405 210309
rect 294095 192309 294111 192587
rect 294389 192309 294405 192587
rect 294095 174587 294405 192309
rect 294095 174309 294111 174587
rect 294389 174309 294405 174587
rect 294095 156587 294405 174309
rect 294095 156309 294111 156587
rect 294389 156309 294405 156587
rect 294095 138587 294405 156309
rect 294095 138309 294111 138587
rect 294389 138309 294405 138587
rect 294095 120587 294405 138309
rect 294095 120309 294111 120587
rect 294389 120309 294405 120587
rect 294095 102587 294405 120309
rect 294095 102309 294111 102587
rect 294389 102309 294405 102587
rect 294095 84587 294405 102309
rect 294095 84309 294111 84587
rect 294389 84309 294405 84587
rect 294095 66587 294405 84309
rect 294095 66309 294111 66587
rect 294389 66309 294405 66587
rect 294095 48587 294405 66309
rect 294095 48309 294111 48587
rect 294389 48309 294405 48587
rect 294095 30587 294405 48309
rect 294095 30309 294111 30587
rect 294389 30309 294405 30587
rect 294095 12587 294405 30309
rect 294095 12309 294111 12587
rect 294389 12309 294405 12587
rect 294095 -1613 294405 12309
rect 294095 -1891 294111 -1613
rect 294389 -1891 294405 -1613
rect 294095 -1907 294405 -1891
rect 294575 347447 294885 354061
rect 294575 347169 294591 347447
rect 294869 347169 294885 347447
rect 294575 329447 294885 347169
rect 294575 329169 294591 329447
rect 294869 329169 294885 329447
rect 294575 311447 294885 329169
rect 294575 311169 294591 311447
rect 294869 311169 294885 311447
rect 294575 293447 294885 311169
rect 294575 293169 294591 293447
rect 294869 293169 294885 293447
rect 294575 275447 294885 293169
rect 294575 275169 294591 275447
rect 294869 275169 294885 275447
rect 294575 257447 294885 275169
rect 294575 257169 294591 257447
rect 294869 257169 294885 257447
rect 294575 239447 294885 257169
rect 294575 239169 294591 239447
rect 294869 239169 294885 239447
rect 294575 221447 294885 239169
rect 294575 221169 294591 221447
rect 294869 221169 294885 221447
rect 294575 203447 294885 221169
rect 294575 203169 294591 203447
rect 294869 203169 294885 203447
rect 294575 185447 294885 203169
rect 294575 185169 294591 185447
rect 294869 185169 294885 185447
rect 294575 167447 294885 185169
rect 294575 167169 294591 167447
rect 294869 167169 294885 167447
rect 294575 149447 294885 167169
rect 294575 149169 294591 149447
rect 294869 149169 294885 149447
rect 294575 131447 294885 149169
rect 294575 131169 294591 131447
rect 294869 131169 294885 131447
rect 294575 113447 294885 131169
rect 294575 113169 294591 113447
rect 294869 113169 294885 113447
rect 294575 95447 294885 113169
rect 294575 95169 294591 95447
rect 294869 95169 294885 95447
rect 294575 77447 294885 95169
rect 294575 77169 294591 77447
rect 294869 77169 294885 77447
rect 294575 59447 294885 77169
rect 294575 59169 294591 59447
rect 294869 59169 294885 59447
rect 294575 41447 294885 59169
rect 294575 41169 294591 41447
rect 294869 41169 294885 41447
rect 294575 23447 294885 41169
rect 294575 23169 294591 23447
rect 294869 23169 294885 23447
rect 294575 5447 294885 23169
rect 294575 5169 294591 5447
rect 294869 5169 294885 5447
rect 294575 -2093 294885 5169
rect 294575 -2371 294591 -2093
rect 294869 -2371 294885 -2093
rect 294575 -2387 294885 -2371
rect 295055 338447 295365 354541
rect 295055 338169 295071 338447
rect 295349 338169 295365 338447
rect 295055 320447 295365 338169
rect 295055 320169 295071 320447
rect 295349 320169 295365 320447
rect 295055 302447 295365 320169
rect 295055 302169 295071 302447
rect 295349 302169 295365 302447
rect 295055 284447 295365 302169
rect 295055 284169 295071 284447
rect 295349 284169 295365 284447
rect 295055 266447 295365 284169
rect 295055 266169 295071 266447
rect 295349 266169 295365 266447
rect 295055 248447 295365 266169
rect 295055 248169 295071 248447
rect 295349 248169 295365 248447
rect 295055 230447 295365 248169
rect 295055 230169 295071 230447
rect 295349 230169 295365 230447
rect 295055 212447 295365 230169
rect 295055 212169 295071 212447
rect 295349 212169 295365 212447
rect 295055 194447 295365 212169
rect 295055 194169 295071 194447
rect 295349 194169 295365 194447
rect 295055 176447 295365 194169
rect 295055 176169 295071 176447
rect 295349 176169 295365 176447
rect 295055 158447 295365 176169
rect 295055 158169 295071 158447
rect 295349 158169 295365 158447
rect 295055 140447 295365 158169
rect 295055 140169 295071 140447
rect 295349 140169 295365 140447
rect 295055 122447 295365 140169
rect 295055 122169 295071 122447
rect 295349 122169 295365 122447
rect 295055 104447 295365 122169
rect 295055 104169 295071 104447
rect 295349 104169 295365 104447
rect 295055 86447 295365 104169
rect 295055 86169 295071 86447
rect 295349 86169 295365 86447
rect 295055 68447 295365 86169
rect 295055 68169 295071 68447
rect 295349 68169 295365 68447
rect 295055 50447 295365 68169
rect 295055 50169 295071 50447
rect 295349 50169 295365 50447
rect 295055 32447 295365 50169
rect 295055 32169 295071 32447
rect 295349 32169 295365 32447
rect 295055 14447 295365 32169
rect 295055 14169 295071 14447
rect 295349 14169 295365 14447
rect 295055 -2573 295365 14169
rect 295055 -2851 295071 -2573
rect 295349 -2851 295365 -2573
rect 295055 -2867 295365 -2851
rect 295535 349307 295845 355021
rect 295535 349029 295551 349307
rect 295829 349029 295845 349307
rect 295535 331307 295845 349029
rect 295535 331029 295551 331307
rect 295829 331029 295845 331307
rect 295535 313307 295845 331029
rect 295535 313029 295551 313307
rect 295829 313029 295845 313307
rect 295535 295307 295845 313029
rect 295535 295029 295551 295307
rect 295829 295029 295845 295307
rect 295535 277307 295845 295029
rect 295535 277029 295551 277307
rect 295829 277029 295845 277307
rect 295535 259307 295845 277029
rect 295535 259029 295551 259307
rect 295829 259029 295845 259307
rect 295535 241307 295845 259029
rect 295535 241029 295551 241307
rect 295829 241029 295845 241307
rect 295535 223307 295845 241029
rect 295535 223029 295551 223307
rect 295829 223029 295845 223307
rect 295535 205307 295845 223029
rect 295535 205029 295551 205307
rect 295829 205029 295845 205307
rect 295535 187307 295845 205029
rect 295535 187029 295551 187307
rect 295829 187029 295845 187307
rect 295535 169307 295845 187029
rect 295535 169029 295551 169307
rect 295829 169029 295845 169307
rect 295535 151307 295845 169029
rect 295535 151029 295551 151307
rect 295829 151029 295845 151307
rect 295535 133307 295845 151029
rect 295535 133029 295551 133307
rect 295829 133029 295845 133307
rect 295535 115307 295845 133029
rect 295535 115029 295551 115307
rect 295829 115029 295845 115307
rect 295535 97307 295845 115029
rect 295535 97029 295551 97307
rect 295829 97029 295845 97307
rect 295535 79307 295845 97029
rect 295535 79029 295551 79307
rect 295829 79029 295845 79307
rect 295535 61307 295845 79029
rect 295535 61029 295551 61307
rect 295829 61029 295845 61307
rect 295535 43307 295845 61029
rect 295535 43029 295551 43307
rect 295829 43029 295845 43307
rect 295535 25307 295845 43029
rect 295535 25029 295551 25307
rect 295829 25029 295845 25307
rect 295535 7307 295845 25029
rect 295535 7029 295551 7307
rect 295829 7029 295845 7307
rect 295535 -3053 295845 7029
rect 295535 -3331 295551 -3053
rect 295829 -3331 295845 -3053
rect 295535 -3347 295845 -3331
rect 296015 340307 296325 355501
rect 296015 340029 296031 340307
rect 296309 340029 296325 340307
rect 296015 322307 296325 340029
rect 296015 322029 296031 322307
rect 296309 322029 296325 322307
rect 296015 304307 296325 322029
rect 296015 304029 296031 304307
rect 296309 304029 296325 304307
rect 296015 286307 296325 304029
rect 296015 286029 296031 286307
rect 296309 286029 296325 286307
rect 296015 268307 296325 286029
rect 296015 268029 296031 268307
rect 296309 268029 296325 268307
rect 296015 250307 296325 268029
rect 296015 250029 296031 250307
rect 296309 250029 296325 250307
rect 296015 232307 296325 250029
rect 296015 232029 296031 232307
rect 296309 232029 296325 232307
rect 296015 214307 296325 232029
rect 296015 214029 296031 214307
rect 296309 214029 296325 214307
rect 296015 196307 296325 214029
rect 296015 196029 296031 196307
rect 296309 196029 296325 196307
rect 296015 178307 296325 196029
rect 296015 178029 296031 178307
rect 296309 178029 296325 178307
rect 296015 160307 296325 178029
rect 296015 160029 296031 160307
rect 296309 160029 296325 160307
rect 296015 142307 296325 160029
rect 296015 142029 296031 142307
rect 296309 142029 296325 142307
rect 296015 124307 296325 142029
rect 296015 124029 296031 124307
rect 296309 124029 296325 124307
rect 296015 106307 296325 124029
rect 296015 106029 296031 106307
rect 296309 106029 296325 106307
rect 296015 88307 296325 106029
rect 296015 88029 296031 88307
rect 296309 88029 296325 88307
rect 296015 70307 296325 88029
rect 296015 70029 296031 70307
rect 296309 70029 296325 70307
rect 296015 52307 296325 70029
rect 296015 52029 296031 52307
rect 296309 52029 296325 52307
rect 296015 34307 296325 52029
rect 296015 34029 296031 34307
rect 296309 34029 296325 34307
rect 296015 16307 296325 34029
rect 296015 16029 296031 16307
rect 296309 16029 296325 16307
rect 285477 -3811 285493 -3533
rect 285771 -3811 285787 -3533
rect 285477 -3827 285787 -3811
rect 296015 -3533 296325 16029
rect 296015 -3811 296031 -3533
rect 296309 -3811 296325 -3533
rect 296015 -3827 296325 -3811
<< via4 >>
rect -4347 355501 -4069 355779
rect -4347 340029 -4069 340307
rect -4347 322029 -4069 322307
rect -4347 304029 -4069 304307
rect -4347 286029 -4069 286307
rect -4347 268029 -4069 268307
rect -4347 250029 -4069 250307
rect -4347 232029 -4069 232307
rect -4347 214029 -4069 214307
rect -4347 196029 -4069 196307
rect -4347 178029 -4069 178307
rect -4347 160029 -4069 160307
rect -4347 142029 -4069 142307
rect -4347 124029 -4069 124307
rect -4347 106029 -4069 106307
rect -4347 88029 -4069 88307
rect -4347 70029 -4069 70307
rect -4347 52029 -4069 52307
rect -4347 34029 -4069 34307
rect -4347 16029 -4069 16307
rect -3867 355021 -3589 355299
rect 6493 355021 6771 355299
rect -3867 349029 -3589 349307
rect -3867 331029 -3589 331307
rect -3867 313029 -3589 313307
rect -3867 295029 -3589 295307
rect -3867 277029 -3589 277307
rect -3867 259029 -3589 259307
rect -3867 241029 -3589 241307
rect -3867 223029 -3589 223307
rect -3867 205029 -3589 205307
rect -3867 187029 -3589 187307
rect -3867 169029 -3589 169307
rect -3867 151029 -3589 151307
rect -3867 133029 -3589 133307
rect -3867 115029 -3589 115307
rect -3867 97029 -3589 97307
rect -3867 79029 -3589 79307
rect -3867 61029 -3589 61307
rect -3867 43029 -3589 43307
rect -3867 25029 -3589 25307
rect -3867 7029 -3589 7307
rect -3387 354541 -3109 354819
rect -3387 338169 -3109 338447
rect -3387 320169 -3109 320447
rect -3387 302169 -3109 302447
rect -3387 284169 -3109 284447
rect -3387 266169 -3109 266447
rect -3387 248169 -3109 248447
rect -3387 230169 -3109 230447
rect -3387 212169 -3109 212447
rect -3387 194169 -3109 194447
rect -3387 176169 -3109 176447
rect -3387 158169 -3109 158447
rect -3387 140169 -3109 140447
rect -3387 122169 -3109 122447
rect -3387 104169 -3109 104447
rect -3387 86169 -3109 86447
rect -3387 68169 -3109 68447
rect -3387 50169 -3109 50447
rect -3387 32169 -3109 32447
rect -3387 14169 -3109 14447
rect -2907 354061 -2629 354339
rect 4633 354061 4911 354339
rect -2907 347169 -2629 347447
rect -2907 329169 -2629 329447
rect -2907 311169 -2629 311447
rect -2907 293169 -2629 293447
rect -2907 275169 -2629 275447
rect -2907 257169 -2629 257447
rect -2907 239169 -2629 239447
rect -2907 221169 -2629 221447
rect -2907 203169 -2629 203447
rect -2907 185169 -2629 185447
rect -2907 167169 -2629 167447
rect -2907 149169 -2629 149447
rect -2907 131169 -2629 131447
rect -2907 113169 -2629 113447
rect -2907 95169 -2629 95447
rect -2907 77169 -2629 77447
rect -2907 59169 -2629 59447
rect -2907 41169 -2629 41447
rect -2907 23169 -2629 23447
rect -2907 5169 -2629 5447
rect -2427 353581 -2149 353859
rect -2427 336309 -2149 336587
rect -2427 318309 -2149 318587
rect -2427 300309 -2149 300587
rect -2427 282309 -2149 282587
rect -2427 264309 -2149 264587
rect -2427 246309 -2149 246587
rect -2427 228309 -2149 228587
rect -2427 210309 -2149 210587
rect -2427 192309 -2149 192587
rect -2427 174309 -2149 174587
rect -2427 156309 -2149 156587
rect -2427 138309 -2149 138587
rect -2427 120309 -2149 120587
rect -2427 102309 -2149 102587
rect -2427 84309 -2149 84587
rect -2427 66309 -2149 66587
rect -2427 48309 -2149 48587
rect -2427 30309 -2149 30587
rect -2427 12309 -2149 12587
rect -1947 353101 -1669 353379
rect 2773 353101 3051 353379
rect -1947 345309 -1669 345587
rect -1947 327309 -1669 327587
rect -1947 309309 -1669 309587
rect -1947 291309 -1669 291587
rect -1947 273309 -1669 273587
rect -1947 255309 -1669 255587
rect -1947 237309 -1669 237587
rect -1947 219309 -1669 219587
rect -1947 201309 -1669 201587
rect -1947 183309 -1669 183587
rect -1947 165309 -1669 165587
rect -1947 147309 -1669 147587
rect -1947 129309 -1669 129587
rect -1947 111309 -1669 111587
rect -1947 93309 -1669 93587
rect -1947 75309 -1669 75587
rect -1947 57309 -1669 57587
rect -1947 39309 -1669 39587
rect -1947 21309 -1669 21587
rect -1947 3309 -1669 3587
rect -1467 352621 -1189 352899
rect -1467 334449 -1189 334727
rect -1467 316449 -1189 316727
rect -1467 298449 -1189 298727
rect -1467 280449 -1189 280727
rect -1467 262449 -1189 262727
rect -1467 244449 -1189 244727
rect -1467 226449 -1189 226727
rect -1467 208449 -1189 208727
rect -1467 190449 -1189 190727
rect -1467 172449 -1189 172727
rect -1467 154449 -1189 154727
rect -1467 136449 -1189 136727
rect -1467 118449 -1189 118727
rect -1467 100449 -1189 100727
rect -1467 82449 -1189 82727
rect -1467 64449 -1189 64727
rect -1467 46449 -1189 46727
rect -1467 28449 -1189 28727
rect -1467 10449 -1189 10727
rect -987 352141 -709 352419
rect -987 343449 -709 343727
rect -987 325449 -709 325727
rect -987 307449 -709 307727
rect -987 289449 -709 289727
rect -987 271449 -709 271727
rect -987 253449 -709 253727
rect -987 235449 -709 235727
rect -987 217449 -709 217727
rect -987 199449 -709 199727
rect -987 181449 -709 181727
rect -987 163449 -709 163727
rect -987 145449 -709 145727
rect -987 127449 -709 127727
rect -987 109449 -709 109727
rect -987 91449 -709 91727
rect -987 73449 -709 73727
rect -987 55449 -709 55727
rect -987 37449 -709 37727
rect -987 19449 -709 19727
rect -987 1449 -709 1727
rect -987 -451 -709 -173
rect 913 352141 1191 352419
rect 913 343449 1191 343727
rect 913 325449 1191 325727
rect 913 307449 1191 307727
rect 913 289449 1191 289727
rect 913 271449 1191 271727
rect 913 253449 1191 253727
rect 913 235449 1191 235727
rect 913 217449 1191 217727
rect 913 199449 1191 199727
rect 913 181449 1191 181727
rect 913 163449 1191 163727
rect 913 145449 1191 145727
rect 913 127449 1191 127727
rect 913 109449 1191 109727
rect 913 91449 1191 91727
rect 913 73449 1191 73727
rect 913 55449 1191 55727
rect 913 37449 1191 37727
rect 913 19449 1191 19727
rect 913 1449 1191 1727
rect 913 -451 1191 -173
rect -1467 -931 -1189 -653
rect 2773 345309 3051 345587
rect 2773 327309 3051 327587
rect 2773 309309 3051 309587
rect 2773 291309 3051 291587
rect 2773 273309 3051 273587
rect 2773 255309 3051 255587
rect 2773 237309 3051 237587
rect 2773 219309 3051 219587
rect 2773 201309 3051 201587
rect 2773 183309 3051 183587
rect 2773 165309 3051 165587
rect 2773 147309 3051 147587
rect 2773 129309 3051 129587
rect 2773 111309 3051 111587
rect 2773 93309 3051 93587
rect 2773 75309 3051 75587
rect 2773 57309 3051 57587
rect 2773 39309 3051 39587
rect 2773 21309 3051 21587
rect 2773 3309 3051 3587
rect -1947 -1411 -1669 -1133
rect 2773 -1411 3051 -1133
rect -2427 -1891 -2149 -1613
rect 4633 347169 4911 347447
rect 4633 329169 4911 329447
rect 4633 311169 4911 311447
rect 4633 293169 4911 293447
rect 4633 275169 4911 275447
rect 4633 257169 4911 257447
rect 4633 239169 4911 239447
rect 4633 221169 4911 221447
rect 4633 203169 4911 203447
rect 4633 185169 4911 185447
rect 4633 167169 4911 167447
rect 4633 149169 4911 149447
rect 4633 131169 4911 131447
rect 4633 113169 4911 113447
rect 4633 95169 4911 95447
rect 4633 77169 4911 77447
rect 4633 59169 4911 59447
rect 4633 41169 4911 41447
rect 4633 23169 4911 23447
rect 4633 5169 4911 5447
rect -2907 -2371 -2629 -2093
rect 4633 -2371 4911 -2093
rect -3387 -2851 -3109 -2573
rect 15493 355501 15771 355779
rect 13633 354541 13911 354819
rect 11773 353581 12051 353859
rect 6493 349029 6771 349307
rect 6493 331029 6771 331307
rect 6493 313029 6771 313307
rect 6493 295029 6771 295307
rect 6493 277029 6771 277307
rect 6493 259029 6771 259307
rect 6493 241029 6771 241307
rect 6493 223029 6771 223307
rect 6493 205029 6771 205307
rect 6493 187029 6771 187307
rect 6493 169029 6771 169307
rect 6493 151029 6771 151307
rect 6493 133029 6771 133307
rect 6493 115029 6771 115307
rect 6493 97029 6771 97307
rect 6493 79029 6771 79307
rect 6493 61029 6771 61307
rect 6493 43029 6771 43307
rect 6493 25029 6771 25307
rect 6493 7029 6771 7307
rect -3867 -3331 -3589 -3053
rect 9913 352621 10191 352899
rect 9913 334449 10191 334727
rect 9913 316449 10191 316727
rect 9913 298449 10191 298727
rect 9913 280449 10191 280727
rect 9913 262449 10191 262727
rect 9913 244449 10191 244727
rect 9913 226449 10191 226727
rect 9913 208449 10191 208727
rect 9913 190449 10191 190727
rect 9913 172449 10191 172727
rect 9913 154449 10191 154727
rect 9913 136449 10191 136727
rect 9913 118449 10191 118727
rect 9913 100449 10191 100727
rect 9913 82449 10191 82727
rect 9913 64449 10191 64727
rect 9913 46449 10191 46727
rect 9913 28449 10191 28727
rect 9913 10449 10191 10727
rect 9913 -931 10191 -653
rect 11773 336309 12051 336587
rect 11773 318309 12051 318587
rect 11773 300309 12051 300587
rect 11773 282309 12051 282587
rect 11773 264309 12051 264587
rect 11773 246309 12051 246587
rect 11773 228309 12051 228587
rect 11773 210309 12051 210587
rect 11773 192309 12051 192587
rect 11773 174309 12051 174587
rect 11773 156309 12051 156587
rect 11773 138309 12051 138587
rect 11773 120309 12051 120587
rect 11773 102309 12051 102587
rect 11773 84309 12051 84587
rect 11773 66309 12051 66587
rect 11773 48309 12051 48587
rect 11773 30309 12051 30587
rect 11773 12309 12051 12587
rect 11773 -1891 12051 -1613
rect 13633 338169 13911 338447
rect 13633 320169 13911 320447
rect 13633 302169 13911 302447
rect 13633 284169 13911 284447
rect 13633 266169 13911 266447
rect 13633 248169 13911 248447
rect 13633 230169 13911 230447
rect 13633 212169 13911 212447
rect 13633 194169 13911 194447
rect 13633 176169 13911 176447
rect 13633 158169 13911 158447
rect 13633 140169 13911 140447
rect 13633 122169 13911 122447
rect 13633 104169 13911 104447
rect 13633 86169 13911 86447
rect 13633 68169 13911 68447
rect 13633 50169 13911 50447
rect 13633 32169 13911 32447
rect 13633 14169 13911 14447
rect 13633 -2851 13911 -2573
rect 24493 355021 24771 355299
rect 22633 354061 22911 354339
rect 20773 353101 21051 353379
rect 15493 340029 15771 340307
rect 15493 322029 15771 322307
rect 15493 304029 15771 304307
rect 15493 286029 15771 286307
rect 15493 268029 15771 268307
rect 15493 250029 15771 250307
rect 15493 232029 15771 232307
rect 15493 214029 15771 214307
rect 15493 196029 15771 196307
rect 15493 178029 15771 178307
rect 15493 160029 15771 160307
rect 15493 142029 15771 142307
rect 15493 124029 15771 124307
rect 15493 106029 15771 106307
rect 15493 88029 15771 88307
rect 15493 70029 15771 70307
rect 15493 52029 15771 52307
rect 15493 34029 15771 34307
rect 15493 16029 15771 16307
rect 6493 -3331 6771 -3053
rect -4347 -3811 -4069 -3533
rect 18913 352141 19191 352419
rect 18913 343449 19191 343727
rect 18913 325449 19191 325727
rect 18913 307449 19191 307727
rect 18913 289449 19191 289727
rect 18913 271449 19191 271727
rect 18913 253449 19191 253727
rect 18913 235449 19191 235727
rect 18913 217449 19191 217727
rect 18913 199449 19191 199727
rect 18913 181449 19191 181727
rect 18913 163449 19191 163727
rect 18913 145449 19191 145727
rect 18913 127449 19191 127727
rect 18913 109449 19191 109727
rect 18913 91449 19191 91727
rect 18913 73449 19191 73727
rect 18913 55449 19191 55727
rect 18913 37449 19191 37727
rect 18913 19449 19191 19727
rect 18913 1449 19191 1727
rect 18913 -451 19191 -173
rect 20773 345309 21051 345587
rect 20773 327309 21051 327587
rect 20773 309309 21051 309587
rect 20773 291309 21051 291587
rect 20773 273309 21051 273587
rect 20773 255309 21051 255587
rect 20773 237309 21051 237587
rect 20773 219309 21051 219587
rect 20773 201309 21051 201587
rect 20773 183309 21051 183587
rect 20773 165309 21051 165587
rect 20773 147309 21051 147587
rect 20773 129309 21051 129587
rect 20773 111309 21051 111587
rect 20773 93309 21051 93587
rect 20773 75309 21051 75587
rect 20773 57309 21051 57587
rect 20773 39309 21051 39587
rect 20773 21309 21051 21587
rect 20773 3309 21051 3587
rect 20773 -1411 21051 -1133
rect 22633 347169 22911 347447
rect 22633 329169 22911 329447
rect 22633 311169 22911 311447
rect 22633 293169 22911 293447
rect 22633 275169 22911 275447
rect 22633 257169 22911 257447
rect 22633 239169 22911 239447
rect 22633 221169 22911 221447
rect 22633 203169 22911 203447
rect 22633 185169 22911 185447
rect 22633 167169 22911 167447
rect 22633 149169 22911 149447
rect 22633 131169 22911 131447
rect 22633 113169 22911 113447
rect 22633 95169 22911 95447
rect 22633 77169 22911 77447
rect 22633 59169 22911 59447
rect 22633 41169 22911 41447
rect 22633 23169 22911 23447
rect 22633 5169 22911 5447
rect 22633 -2371 22911 -2093
rect 33493 355501 33771 355779
rect 31633 354541 31911 354819
rect 29773 353581 30051 353859
rect 24493 349029 24771 349307
rect 24493 331029 24771 331307
rect 24493 313029 24771 313307
rect 24493 295029 24771 295307
rect 24493 277029 24771 277307
rect 24493 259029 24771 259307
rect 24493 241029 24771 241307
rect 24493 223029 24771 223307
rect 24493 205029 24771 205307
rect 24493 187029 24771 187307
rect 24493 169029 24771 169307
rect 24493 151029 24771 151307
rect 24493 133029 24771 133307
rect 24493 115029 24771 115307
rect 24493 97029 24771 97307
rect 24493 79029 24771 79307
rect 24493 61029 24771 61307
rect 24493 43029 24771 43307
rect 24493 25029 24771 25307
rect 24493 7029 24771 7307
rect 15493 -3811 15771 -3533
rect 27913 352621 28191 352899
rect 27913 334449 28191 334727
rect 27913 316449 28191 316727
rect 27913 298449 28191 298727
rect 27913 280449 28191 280727
rect 27913 262449 28191 262727
rect 27913 244449 28191 244727
rect 27913 226449 28191 226727
rect 27913 208449 28191 208727
rect 27913 190449 28191 190727
rect 27913 172449 28191 172727
rect 27913 154449 28191 154727
rect 27913 136449 28191 136727
rect 27913 118449 28191 118727
rect 27913 100449 28191 100727
rect 27913 82449 28191 82727
rect 27913 64449 28191 64727
rect 27913 46449 28191 46727
rect 27913 28449 28191 28727
rect 27913 10449 28191 10727
rect 27913 -931 28191 -653
rect 29773 336309 30051 336587
rect 29773 318309 30051 318587
rect 29773 300309 30051 300587
rect 29773 282309 30051 282587
rect 29773 264309 30051 264587
rect 29773 246309 30051 246587
rect 29773 228309 30051 228587
rect 29773 210309 30051 210587
rect 29773 192309 30051 192587
rect 29773 174309 30051 174587
rect 29773 156309 30051 156587
rect 29773 138309 30051 138587
rect 29773 120309 30051 120587
rect 29773 102309 30051 102587
rect 29773 84309 30051 84587
rect 29773 66309 30051 66587
rect 29773 48309 30051 48587
rect 29773 30309 30051 30587
rect 29773 12309 30051 12587
rect 29773 -1891 30051 -1613
rect 31633 338169 31911 338447
rect 31633 320169 31911 320447
rect 31633 302169 31911 302447
rect 31633 284169 31911 284447
rect 31633 266169 31911 266447
rect 31633 248169 31911 248447
rect 31633 230169 31911 230447
rect 31633 212169 31911 212447
rect 31633 194169 31911 194447
rect 31633 176169 31911 176447
rect 31633 158169 31911 158447
rect 31633 140169 31911 140447
rect 31633 122169 31911 122447
rect 31633 104169 31911 104447
rect 31633 86169 31911 86447
rect 31633 68169 31911 68447
rect 31633 50169 31911 50447
rect 31633 32169 31911 32447
rect 31633 14169 31911 14447
rect 31633 -2851 31911 -2573
rect 42493 355021 42771 355299
rect 40633 354061 40911 354339
rect 38773 353101 39051 353379
rect 33493 340029 33771 340307
rect 33493 322029 33771 322307
rect 33493 304029 33771 304307
rect 33493 286029 33771 286307
rect 33493 268029 33771 268307
rect 33493 250029 33771 250307
rect 33493 232029 33771 232307
rect 33493 214029 33771 214307
rect 33493 196029 33771 196307
rect 33493 178029 33771 178307
rect 33493 160029 33771 160307
rect 33493 142029 33771 142307
rect 33493 124029 33771 124307
rect 33493 106029 33771 106307
rect 33493 88029 33771 88307
rect 33493 70029 33771 70307
rect 33493 52029 33771 52307
rect 33493 34029 33771 34307
rect 33493 16029 33771 16307
rect 24493 -3331 24771 -3053
rect 36913 352141 37191 352419
rect 36913 343449 37191 343727
rect 36913 325449 37191 325727
rect 36913 307449 37191 307727
rect 36913 289449 37191 289727
rect 36913 271449 37191 271727
rect 36913 253449 37191 253727
rect 36913 235449 37191 235727
rect 36913 217449 37191 217727
rect 36913 199449 37191 199727
rect 36913 181449 37191 181727
rect 36913 163449 37191 163727
rect 36913 145449 37191 145727
rect 36913 127449 37191 127727
rect 36913 109449 37191 109727
rect 36913 91449 37191 91727
rect 36913 73449 37191 73727
rect 36913 55449 37191 55727
rect 36913 37449 37191 37727
rect 36913 19449 37191 19727
rect 36913 1449 37191 1727
rect 36913 -451 37191 -173
rect 38773 345309 39051 345587
rect 38773 327309 39051 327587
rect 38773 309309 39051 309587
rect 38773 291309 39051 291587
rect 38773 273309 39051 273587
rect 38773 255309 39051 255587
rect 38773 237309 39051 237587
rect 38773 219309 39051 219587
rect 38773 201309 39051 201587
rect 38773 183309 39051 183587
rect 38773 165309 39051 165587
rect 38773 147309 39051 147587
rect 38773 129309 39051 129587
rect 38773 111309 39051 111587
rect 38773 93309 39051 93587
rect 38773 75309 39051 75587
rect 38773 57309 39051 57587
rect 38773 39309 39051 39587
rect 38773 21309 39051 21587
rect 38773 3309 39051 3587
rect 38773 -1411 39051 -1133
rect 40633 347169 40911 347447
rect 40633 329169 40911 329447
rect 40633 311169 40911 311447
rect 40633 293169 40911 293447
rect 40633 275169 40911 275447
rect 40633 257169 40911 257447
rect 40633 239169 40911 239447
rect 40633 221169 40911 221447
rect 40633 203169 40911 203447
rect 40633 185169 40911 185447
rect 40633 167169 40911 167447
rect 40633 149169 40911 149447
rect 40633 131169 40911 131447
rect 40633 113169 40911 113447
rect 40633 95169 40911 95447
rect 40633 77169 40911 77447
rect 40633 59169 40911 59447
rect 40633 41169 40911 41447
rect 40633 23169 40911 23447
rect 40633 5169 40911 5447
rect 40633 -2371 40911 -2093
rect 51493 355501 51771 355779
rect 49633 354541 49911 354819
rect 47773 353581 48051 353859
rect 42493 349029 42771 349307
rect 42493 331029 42771 331307
rect 42493 313029 42771 313307
rect 42493 295029 42771 295307
rect 42493 277029 42771 277307
rect 42493 259029 42771 259307
rect 42493 241029 42771 241307
rect 42493 223029 42771 223307
rect 42493 205029 42771 205307
rect 42493 187029 42771 187307
rect 42493 169029 42771 169307
rect 42493 151029 42771 151307
rect 42493 133029 42771 133307
rect 42493 115029 42771 115307
rect 42493 97029 42771 97307
rect 42493 79029 42771 79307
rect 42493 61029 42771 61307
rect 42493 43029 42771 43307
rect 42493 25029 42771 25307
rect 42493 7029 42771 7307
rect 33493 -3811 33771 -3533
rect 45913 352621 46191 352899
rect 45913 334449 46191 334727
rect 45913 316449 46191 316727
rect 45913 298449 46191 298727
rect 45913 280449 46191 280727
rect 45913 262449 46191 262727
rect 45913 244449 46191 244727
rect 45913 226449 46191 226727
rect 45913 208449 46191 208727
rect 45913 190449 46191 190727
rect 45913 172449 46191 172727
rect 45913 154449 46191 154727
rect 45913 136449 46191 136727
rect 45913 118449 46191 118727
rect 45913 100449 46191 100727
rect 45913 82449 46191 82727
rect 45913 64449 46191 64727
rect 45913 46449 46191 46727
rect 45913 28449 46191 28727
rect 45913 10449 46191 10727
rect 45913 -931 46191 -653
rect 47773 336309 48051 336587
rect 47773 318309 48051 318587
rect 47773 300309 48051 300587
rect 47773 282309 48051 282587
rect 47773 264309 48051 264587
rect 47773 246309 48051 246587
rect 47773 228309 48051 228587
rect 47773 210309 48051 210587
rect 47773 192309 48051 192587
rect 47773 174309 48051 174587
rect 47773 156309 48051 156587
rect 47773 138309 48051 138587
rect 47773 120309 48051 120587
rect 47773 102309 48051 102587
rect 47773 84309 48051 84587
rect 47773 66309 48051 66587
rect 47773 48309 48051 48587
rect 47773 30309 48051 30587
rect 47773 12309 48051 12587
rect 47773 -1891 48051 -1613
rect 49633 338169 49911 338447
rect 49633 320169 49911 320447
rect 49633 302169 49911 302447
rect 49633 284169 49911 284447
rect 49633 266169 49911 266447
rect 49633 248169 49911 248447
rect 49633 230169 49911 230447
rect 49633 212169 49911 212447
rect 49633 194169 49911 194447
rect 49633 176169 49911 176447
rect 49633 158169 49911 158447
rect 49633 140169 49911 140447
rect 49633 122169 49911 122447
rect 49633 104169 49911 104447
rect 49633 86169 49911 86447
rect 49633 68169 49911 68447
rect 49633 50169 49911 50447
rect 49633 32169 49911 32447
rect 49633 14169 49911 14447
rect 49633 -2851 49911 -2573
rect 60493 355021 60771 355299
rect 58633 354061 58911 354339
rect 56773 353101 57051 353379
rect 51493 340029 51771 340307
rect 51493 322029 51771 322307
rect 51493 304029 51771 304307
rect 51493 286029 51771 286307
rect 51493 268029 51771 268307
rect 51493 250029 51771 250307
rect 51493 232029 51771 232307
rect 51493 214029 51771 214307
rect 51493 196029 51771 196307
rect 51493 178029 51771 178307
rect 51493 160029 51771 160307
rect 51493 142029 51771 142307
rect 51493 124029 51771 124307
rect 51493 106029 51771 106307
rect 51493 88029 51771 88307
rect 51493 70029 51771 70307
rect 51493 52029 51771 52307
rect 51493 34029 51771 34307
rect 51493 16029 51771 16307
rect 42493 -3331 42771 -3053
rect 54913 352141 55191 352419
rect 54913 343449 55191 343727
rect 54913 325449 55191 325727
rect 54913 307449 55191 307727
rect 54913 289449 55191 289727
rect 54913 271449 55191 271727
rect 54913 253449 55191 253727
rect 54913 235449 55191 235727
rect 54913 217449 55191 217727
rect 54913 199449 55191 199727
rect 54913 181449 55191 181727
rect 54913 163449 55191 163727
rect 54913 145449 55191 145727
rect 54913 127449 55191 127727
rect 54913 109449 55191 109727
rect 54913 91449 55191 91727
rect 54913 73449 55191 73727
rect 54913 55449 55191 55727
rect 54913 37449 55191 37727
rect 54913 19449 55191 19727
rect 54913 1449 55191 1727
rect 54913 -451 55191 -173
rect 56773 345309 57051 345587
rect 56773 327309 57051 327587
rect 56773 309309 57051 309587
rect 56773 291309 57051 291587
rect 56773 273309 57051 273587
rect 56773 255309 57051 255587
rect 56773 237309 57051 237587
rect 56773 219309 57051 219587
rect 56773 201309 57051 201587
rect 56773 183309 57051 183587
rect 56773 165309 57051 165587
rect 56773 147309 57051 147587
rect 56773 129309 57051 129587
rect 56773 111309 57051 111587
rect 56773 93309 57051 93587
rect 56773 75309 57051 75587
rect 56773 57309 57051 57587
rect 56773 39309 57051 39587
rect 56773 21309 57051 21587
rect 56773 3309 57051 3587
rect 56773 -1411 57051 -1133
rect 58633 347169 58911 347447
rect 58633 329169 58911 329447
rect 58633 311169 58911 311447
rect 58633 293169 58911 293447
rect 58633 275169 58911 275447
rect 58633 257169 58911 257447
rect 58633 239169 58911 239447
rect 58633 221169 58911 221447
rect 58633 203169 58911 203447
rect 58633 185169 58911 185447
rect 58633 167169 58911 167447
rect 58633 149169 58911 149447
rect 58633 131169 58911 131447
rect 58633 113169 58911 113447
rect 58633 95169 58911 95447
rect 58633 77169 58911 77447
rect 58633 59169 58911 59447
rect 58633 41169 58911 41447
rect 58633 23169 58911 23447
rect 58633 5169 58911 5447
rect 58633 -2371 58911 -2093
rect 69493 355501 69771 355779
rect 67633 354541 67911 354819
rect 65773 353581 66051 353859
rect 60493 349029 60771 349307
rect 60493 331029 60771 331307
rect 60493 313029 60771 313307
rect 60493 295029 60771 295307
rect 60493 277029 60771 277307
rect 60493 259029 60771 259307
rect 60493 241029 60771 241307
rect 60493 223029 60771 223307
rect 60493 205029 60771 205307
rect 60493 187029 60771 187307
rect 60493 169029 60771 169307
rect 60493 151029 60771 151307
rect 60493 133029 60771 133307
rect 60493 115029 60771 115307
rect 60493 97029 60771 97307
rect 60493 79029 60771 79307
rect 60493 61029 60771 61307
rect 60493 43029 60771 43307
rect 60493 25029 60771 25307
rect 60493 7029 60771 7307
rect 51493 -3811 51771 -3533
rect 63913 352621 64191 352899
rect 63913 334449 64191 334727
rect 63913 316449 64191 316727
rect 63913 298449 64191 298727
rect 63913 280449 64191 280727
rect 63913 262449 64191 262727
rect 63913 244449 64191 244727
rect 63913 226449 64191 226727
rect 63913 208449 64191 208727
rect 63913 190449 64191 190727
rect 63913 172449 64191 172727
rect 63913 154449 64191 154727
rect 63913 136449 64191 136727
rect 63913 118449 64191 118727
rect 63913 100449 64191 100727
rect 63913 82449 64191 82727
rect 63913 64449 64191 64727
rect 63913 46449 64191 46727
rect 63913 28449 64191 28727
rect 63913 10449 64191 10727
rect 63913 -931 64191 -653
rect 65773 336309 66051 336587
rect 65773 318309 66051 318587
rect 65773 300309 66051 300587
rect 65773 282309 66051 282587
rect 65773 264309 66051 264587
rect 65773 246309 66051 246587
rect 65773 228309 66051 228587
rect 65773 210309 66051 210587
rect 65773 192309 66051 192587
rect 65773 174309 66051 174587
rect 65773 156309 66051 156587
rect 65773 138309 66051 138587
rect 65773 120309 66051 120587
rect 65773 102309 66051 102587
rect 65773 84309 66051 84587
rect 65773 66309 66051 66587
rect 65773 48309 66051 48587
rect 65773 30309 66051 30587
rect 65773 12309 66051 12587
rect 65773 -1891 66051 -1613
rect 67633 338169 67911 338447
rect 67633 320169 67911 320447
rect 67633 302169 67911 302447
rect 67633 284169 67911 284447
rect 67633 266169 67911 266447
rect 67633 248169 67911 248447
rect 67633 230169 67911 230447
rect 67633 212169 67911 212447
rect 67633 194169 67911 194447
rect 67633 176169 67911 176447
rect 67633 158169 67911 158447
rect 67633 140169 67911 140447
rect 67633 122169 67911 122447
rect 67633 104169 67911 104447
rect 67633 86169 67911 86447
rect 67633 68169 67911 68447
rect 67633 50169 67911 50447
rect 67633 32169 67911 32447
rect 67633 14169 67911 14447
rect 67633 -2851 67911 -2573
rect 78493 355021 78771 355299
rect 76633 354061 76911 354339
rect 74773 353101 75051 353379
rect 69493 340029 69771 340307
rect 69493 322029 69771 322307
rect 69493 304029 69771 304307
rect 69493 286029 69771 286307
rect 69493 268029 69771 268307
rect 69493 250029 69771 250307
rect 69493 232029 69771 232307
rect 69493 214029 69771 214307
rect 69493 196029 69771 196307
rect 69493 178029 69771 178307
rect 69493 160029 69771 160307
rect 69493 142029 69771 142307
rect 69493 124029 69771 124307
rect 69493 106029 69771 106307
rect 69493 88029 69771 88307
rect 69493 70029 69771 70307
rect 69493 52029 69771 52307
rect 69493 34029 69771 34307
rect 69493 16029 69771 16307
rect 60493 -3331 60771 -3053
rect 72913 352141 73191 352419
rect 72913 343449 73191 343727
rect 72913 325449 73191 325727
rect 72913 307449 73191 307727
rect 72913 289449 73191 289727
rect 72913 271449 73191 271727
rect 72913 253449 73191 253727
rect 72913 235449 73191 235727
rect 72913 217449 73191 217727
rect 72913 199449 73191 199727
rect 72913 181449 73191 181727
rect 72913 163449 73191 163727
rect 72913 145449 73191 145727
rect 72913 127449 73191 127727
rect 72913 109449 73191 109727
rect 72913 91449 73191 91727
rect 72913 73449 73191 73727
rect 72913 55449 73191 55727
rect 72913 37449 73191 37727
rect 72913 19449 73191 19727
rect 72913 1449 73191 1727
rect 72913 -451 73191 -173
rect 74773 345309 75051 345587
rect 74773 327309 75051 327587
rect 74773 309309 75051 309587
rect 74773 291309 75051 291587
rect 74773 273309 75051 273587
rect 74773 255309 75051 255587
rect 74773 237309 75051 237587
rect 74773 219309 75051 219587
rect 74773 201309 75051 201587
rect 74773 183309 75051 183587
rect 74773 165309 75051 165587
rect 74773 147309 75051 147587
rect 74773 129309 75051 129587
rect 74773 111309 75051 111587
rect 74773 93309 75051 93587
rect 74773 75309 75051 75587
rect 74773 57309 75051 57587
rect 74773 39309 75051 39587
rect 74773 21309 75051 21587
rect 74773 3309 75051 3587
rect 74773 -1411 75051 -1133
rect 76633 347169 76911 347447
rect 76633 329169 76911 329447
rect 76633 311169 76911 311447
rect 76633 293169 76911 293447
rect 76633 275169 76911 275447
rect 76633 257169 76911 257447
rect 76633 239169 76911 239447
rect 76633 221169 76911 221447
rect 76633 203169 76911 203447
rect 76633 185169 76911 185447
rect 76633 167169 76911 167447
rect 76633 149169 76911 149447
rect 76633 131169 76911 131447
rect 76633 113169 76911 113447
rect 76633 95169 76911 95447
rect 76633 77169 76911 77447
rect 76633 59169 76911 59447
rect 76633 41169 76911 41447
rect 76633 23169 76911 23447
rect 76633 5169 76911 5447
rect 76633 -2371 76911 -2093
rect 87493 355501 87771 355779
rect 85633 354541 85911 354819
rect 83773 353581 84051 353859
rect 78493 349029 78771 349307
rect 78493 331029 78771 331307
rect 78493 313029 78771 313307
rect 78493 295029 78771 295307
rect 78493 277029 78771 277307
rect 78493 259029 78771 259307
rect 78493 241029 78771 241307
rect 78493 223029 78771 223307
rect 78493 205029 78771 205307
rect 78493 187029 78771 187307
rect 78493 169029 78771 169307
rect 78493 151029 78771 151307
rect 78493 133029 78771 133307
rect 78493 115029 78771 115307
rect 78493 97029 78771 97307
rect 78493 79029 78771 79307
rect 78493 61029 78771 61307
rect 78493 43029 78771 43307
rect 78493 25029 78771 25307
rect 78493 7029 78771 7307
rect 69493 -3811 69771 -3533
rect 81913 352621 82191 352899
rect 81913 334449 82191 334727
rect 81913 316449 82191 316727
rect 81913 298449 82191 298727
rect 81913 280449 82191 280727
rect 81913 262449 82191 262727
rect 81913 244449 82191 244727
rect 81913 226449 82191 226727
rect 81913 208449 82191 208727
rect 81913 190449 82191 190727
rect 81913 172449 82191 172727
rect 81913 154449 82191 154727
rect 81913 136449 82191 136727
rect 81913 118449 82191 118727
rect 81913 100449 82191 100727
rect 81913 82449 82191 82727
rect 81913 64449 82191 64727
rect 81913 46449 82191 46727
rect 81913 28449 82191 28727
rect 81913 10449 82191 10727
rect 81913 -931 82191 -653
rect 83773 336309 84051 336587
rect 83773 318309 84051 318587
rect 83773 300309 84051 300587
rect 83773 282309 84051 282587
rect 83773 264309 84051 264587
rect 83773 246309 84051 246587
rect 83773 228309 84051 228587
rect 83773 210309 84051 210587
rect 83773 192309 84051 192587
rect 83773 174309 84051 174587
rect 83773 156309 84051 156587
rect 83773 138309 84051 138587
rect 83773 120309 84051 120587
rect 83773 102309 84051 102587
rect 83773 84309 84051 84587
rect 83773 66309 84051 66587
rect 83773 48309 84051 48587
rect 83773 30309 84051 30587
rect 83773 12309 84051 12587
rect 83773 -1891 84051 -1613
rect 85633 338169 85911 338447
rect 85633 320169 85911 320447
rect 85633 302169 85911 302447
rect 85633 284169 85911 284447
rect 85633 266169 85911 266447
rect 85633 248169 85911 248447
rect 85633 230169 85911 230447
rect 85633 212169 85911 212447
rect 85633 194169 85911 194447
rect 85633 176169 85911 176447
rect 85633 158169 85911 158447
rect 85633 140169 85911 140447
rect 85633 122169 85911 122447
rect 85633 104169 85911 104447
rect 85633 86169 85911 86447
rect 85633 68169 85911 68447
rect 85633 50169 85911 50447
rect 85633 32169 85911 32447
rect 85633 14169 85911 14447
rect 85633 -2851 85911 -2573
rect 96493 355021 96771 355299
rect 94633 354061 94911 354339
rect 92773 353101 93051 353379
rect 87493 340029 87771 340307
rect 87493 322029 87771 322307
rect 87493 304029 87771 304307
rect 87493 286029 87771 286307
rect 87493 268029 87771 268307
rect 87493 250029 87771 250307
rect 87493 232029 87771 232307
rect 87493 214029 87771 214307
rect 87493 196029 87771 196307
rect 87493 178029 87771 178307
rect 87493 160029 87771 160307
rect 87493 142029 87771 142307
rect 87493 124029 87771 124307
rect 87493 106029 87771 106307
rect 87493 88029 87771 88307
rect 87493 70029 87771 70307
rect 87493 52029 87771 52307
rect 87493 34029 87771 34307
rect 87493 16029 87771 16307
rect 78493 -3331 78771 -3053
rect 90913 352141 91191 352419
rect 90913 343449 91191 343727
rect 90913 325449 91191 325727
rect 90913 307449 91191 307727
rect 90913 289449 91191 289727
rect 90913 271449 91191 271727
rect 90913 253449 91191 253727
rect 90913 235449 91191 235727
rect 90913 217449 91191 217727
rect 90913 199449 91191 199727
rect 90913 181449 91191 181727
rect 90913 163449 91191 163727
rect 90913 145449 91191 145727
rect 90913 127449 91191 127727
rect 90913 109449 91191 109727
rect 90913 91449 91191 91727
rect 90913 73449 91191 73727
rect 90913 55449 91191 55727
rect 90913 37449 91191 37727
rect 90913 19449 91191 19727
rect 90913 1449 91191 1727
rect 90913 -451 91191 -173
rect 92773 345309 93051 345587
rect 92773 327309 93051 327587
rect 92773 309309 93051 309587
rect 92773 291309 93051 291587
rect 92773 273309 93051 273587
rect 92773 255309 93051 255587
rect 92773 237309 93051 237587
rect 92773 219309 93051 219587
rect 92773 201309 93051 201587
rect 92773 183309 93051 183587
rect 92773 165309 93051 165587
rect 92773 147309 93051 147587
rect 92773 129309 93051 129587
rect 92773 111309 93051 111587
rect 92773 93309 93051 93587
rect 92773 75309 93051 75587
rect 92773 57309 93051 57587
rect 92773 39309 93051 39587
rect 92773 21309 93051 21587
rect 92773 3309 93051 3587
rect 92773 -1411 93051 -1133
rect 94633 347169 94911 347447
rect 94633 329169 94911 329447
rect 94633 311169 94911 311447
rect 94633 293169 94911 293447
rect 94633 275169 94911 275447
rect 94633 257169 94911 257447
rect 94633 239169 94911 239447
rect 94633 221169 94911 221447
rect 94633 203169 94911 203447
rect 94633 185169 94911 185447
rect 94633 167169 94911 167447
rect 94633 149169 94911 149447
rect 94633 131169 94911 131447
rect 94633 113169 94911 113447
rect 94633 95169 94911 95447
rect 94633 77169 94911 77447
rect 94633 59169 94911 59447
rect 94633 41169 94911 41447
rect 94633 23169 94911 23447
rect 94633 5169 94911 5447
rect 94633 -2371 94911 -2093
rect 105493 355501 105771 355779
rect 103633 354541 103911 354819
rect 101773 353581 102051 353859
rect 96493 349029 96771 349307
rect 96493 331029 96771 331307
rect 96493 313029 96771 313307
rect 96493 295029 96771 295307
rect 96493 277029 96771 277307
rect 96493 259029 96771 259307
rect 96493 241029 96771 241307
rect 96493 223029 96771 223307
rect 96493 205029 96771 205307
rect 96493 187029 96771 187307
rect 96493 169029 96771 169307
rect 96493 151029 96771 151307
rect 96493 133029 96771 133307
rect 96493 115029 96771 115307
rect 96493 97029 96771 97307
rect 96493 79029 96771 79307
rect 96493 61029 96771 61307
rect 96493 43029 96771 43307
rect 96493 25029 96771 25307
rect 96493 7029 96771 7307
rect 87493 -3811 87771 -3533
rect 99913 352621 100191 352899
rect 99913 334449 100191 334727
rect 99913 316449 100191 316727
rect 99913 298449 100191 298727
rect 99913 280449 100191 280727
rect 99913 262449 100191 262727
rect 99913 244449 100191 244727
rect 99913 226449 100191 226727
rect 99913 208449 100191 208727
rect 99913 190449 100191 190727
rect 99913 172449 100191 172727
rect 99913 154449 100191 154727
rect 99913 136449 100191 136727
rect 99913 118449 100191 118727
rect 99913 100449 100191 100727
rect 99913 82449 100191 82727
rect 99913 64449 100191 64727
rect 99913 46449 100191 46727
rect 99913 28449 100191 28727
rect 99913 10449 100191 10727
rect 99913 -931 100191 -653
rect 101773 336309 102051 336587
rect 101773 318309 102051 318587
rect 101773 300309 102051 300587
rect 101773 282309 102051 282587
rect 101773 264309 102051 264587
rect 101773 246309 102051 246587
rect 101773 228309 102051 228587
rect 101773 210309 102051 210587
rect 101773 192309 102051 192587
rect 101773 174309 102051 174587
rect 101773 156309 102051 156587
rect 101773 138309 102051 138587
rect 101773 120309 102051 120587
rect 101773 102309 102051 102587
rect 101773 84309 102051 84587
rect 101773 66309 102051 66587
rect 101773 48309 102051 48587
rect 101773 30309 102051 30587
rect 101773 12309 102051 12587
rect 101773 -1891 102051 -1613
rect 103633 338169 103911 338447
rect 103633 320169 103911 320447
rect 103633 302169 103911 302447
rect 103633 284169 103911 284447
rect 103633 266169 103911 266447
rect 103633 248169 103911 248447
rect 103633 230169 103911 230447
rect 103633 212169 103911 212447
rect 103633 194169 103911 194447
rect 103633 176169 103911 176447
rect 103633 158169 103911 158447
rect 103633 140169 103911 140447
rect 103633 122169 103911 122447
rect 103633 104169 103911 104447
rect 103633 86169 103911 86447
rect 103633 68169 103911 68447
rect 103633 50169 103911 50447
rect 103633 32169 103911 32447
rect 103633 14169 103911 14447
rect 103633 -2851 103911 -2573
rect 114493 355021 114771 355299
rect 112633 354061 112911 354339
rect 110773 353101 111051 353379
rect 105493 340029 105771 340307
rect 105493 322029 105771 322307
rect 105493 304029 105771 304307
rect 105493 286029 105771 286307
rect 105493 268029 105771 268307
rect 105493 250029 105771 250307
rect 105493 232029 105771 232307
rect 105493 214029 105771 214307
rect 105493 196029 105771 196307
rect 105493 178029 105771 178307
rect 105493 160029 105771 160307
rect 105493 142029 105771 142307
rect 105493 124029 105771 124307
rect 105493 106029 105771 106307
rect 105493 88029 105771 88307
rect 105493 70029 105771 70307
rect 105493 52029 105771 52307
rect 105493 34029 105771 34307
rect 105493 16029 105771 16307
rect 96493 -3331 96771 -3053
rect 108913 352141 109191 352419
rect 108913 343449 109191 343727
rect 108913 325449 109191 325727
rect 108913 307449 109191 307727
rect 108913 289449 109191 289727
rect 108913 271449 109191 271727
rect 108913 253449 109191 253727
rect 108913 235449 109191 235727
rect 108913 217449 109191 217727
rect 108913 199449 109191 199727
rect 108913 181449 109191 181727
rect 108913 163449 109191 163727
rect 108913 145449 109191 145727
rect 108913 127449 109191 127727
rect 108913 109449 109191 109727
rect 108913 91449 109191 91727
rect 108913 73449 109191 73727
rect 108913 55449 109191 55727
rect 108913 37449 109191 37727
rect 108913 19449 109191 19727
rect 108913 1449 109191 1727
rect 108913 -451 109191 -173
rect 110773 345309 111051 345587
rect 110773 327309 111051 327587
rect 110773 309309 111051 309587
rect 110773 291309 111051 291587
rect 110773 273309 111051 273587
rect 110773 255309 111051 255587
rect 110773 237309 111051 237587
rect 110773 219309 111051 219587
rect 110773 201309 111051 201587
rect 110773 183309 111051 183587
rect 110773 165309 111051 165587
rect 110773 147309 111051 147587
rect 110773 129309 111051 129587
rect 110773 111309 111051 111587
rect 110773 93309 111051 93587
rect 110773 75309 111051 75587
rect 110773 57309 111051 57587
rect 110773 39309 111051 39587
rect 110773 21309 111051 21587
rect 110773 3309 111051 3587
rect 110773 -1411 111051 -1133
rect 112633 347169 112911 347447
rect 112633 329169 112911 329447
rect 112633 311169 112911 311447
rect 112633 293169 112911 293447
rect 112633 275169 112911 275447
rect 112633 257169 112911 257447
rect 112633 239169 112911 239447
rect 112633 221169 112911 221447
rect 112633 203169 112911 203447
rect 112633 185169 112911 185447
rect 112633 167169 112911 167447
rect 112633 149169 112911 149447
rect 112633 131169 112911 131447
rect 112633 113169 112911 113447
rect 112633 95169 112911 95447
rect 112633 77169 112911 77447
rect 112633 59169 112911 59447
rect 112633 41169 112911 41447
rect 112633 23169 112911 23447
rect 112633 5169 112911 5447
rect 112633 -2371 112911 -2093
rect 123493 355501 123771 355779
rect 121633 354541 121911 354819
rect 119773 353581 120051 353859
rect 114493 349029 114771 349307
rect 114493 331029 114771 331307
rect 114493 313029 114771 313307
rect 114493 295029 114771 295307
rect 114493 277029 114771 277307
rect 114493 259029 114771 259307
rect 114493 241029 114771 241307
rect 114493 223029 114771 223307
rect 114493 205029 114771 205307
rect 114493 187029 114771 187307
rect 114493 169029 114771 169307
rect 114493 151029 114771 151307
rect 114493 133029 114771 133307
rect 114493 115029 114771 115307
rect 114493 97029 114771 97307
rect 114493 79029 114771 79307
rect 114493 61029 114771 61307
rect 114493 43029 114771 43307
rect 114493 25029 114771 25307
rect 114493 7029 114771 7307
rect 105493 -3811 105771 -3533
rect 117913 352621 118191 352899
rect 117913 334449 118191 334727
rect 117913 316449 118191 316727
rect 117913 298449 118191 298727
rect 117913 280449 118191 280727
rect 117913 262449 118191 262727
rect 117913 244449 118191 244727
rect 117913 226449 118191 226727
rect 117913 208449 118191 208727
rect 117913 190449 118191 190727
rect 117913 172449 118191 172727
rect 117913 154449 118191 154727
rect 117913 136449 118191 136727
rect 117913 118449 118191 118727
rect 117913 100449 118191 100727
rect 117913 82449 118191 82727
rect 117913 64449 118191 64727
rect 117913 46449 118191 46727
rect 117913 28449 118191 28727
rect 117913 10449 118191 10727
rect 117913 -931 118191 -653
rect 119773 336309 120051 336587
rect 119773 318309 120051 318587
rect 119773 300309 120051 300587
rect 119773 282309 120051 282587
rect 119773 264309 120051 264587
rect 119773 246309 120051 246587
rect 119773 228309 120051 228587
rect 119773 210309 120051 210587
rect 119773 192309 120051 192587
rect 119773 174309 120051 174587
rect 119773 156309 120051 156587
rect 119773 138309 120051 138587
rect 119773 120309 120051 120587
rect 119773 102309 120051 102587
rect 119773 84309 120051 84587
rect 119773 66309 120051 66587
rect 119773 48309 120051 48587
rect 119773 30309 120051 30587
rect 119773 12309 120051 12587
rect 119773 -1891 120051 -1613
rect 121633 338169 121911 338447
rect 121633 320169 121911 320447
rect 121633 302169 121911 302447
rect 121633 284169 121911 284447
rect 121633 266169 121911 266447
rect 121633 248169 121911 248447
rect 121633 230169 121911 230447
rect 121633 212169 121911 212447
rect 121633 194169 121911 194447
rect 121633 176169 121911 176447
rect 121633 158169 121911 158447
rect 121633 140169 121911 140447
rect 121633 122169 121911 122447
rect 121633 104169 121911 104447
rect 121633 86169 121911 86447
rect 121633 68169 121911 68447
rect 121633 50169 121911 50447
rect 121633 32169 121911 32447
rect 121633 14169 121911 14447
rect 121633 -2851 121911 -2573
rect 132493 355021 132771 355299
rect 130633 354061 130911 354339
rect 128773 353101 129051 353379
rect 123493 340029 123771 340307
rect 123493 322029 123771 322307
rect 123493 304029 123771 304307
rect 123493 286029 123771 286307
rect 123493 268029 123771 268307
rect 123493 250029 123771 250307
rect 123493 232029 123771 232307
rect 123493 214029 123771 214307
rect 123493 196029 123771 196307
rect 123493 178029 123771 178307
rect 123493 160029 123771 160307
rect 123493 142029 123771 142307
rect 123493 124029 123771 124307
rect 123493 106029 123771 106307
rect 123493 88029 123771 88307
rect 123493 70029 123771 70307
rect 123493 52029 123771 52307
rect 123493 34029 123771 34307
rect 123493 16029 123771 16307
rect 114493 -3331 114771 -3053
rect 126913 352141 127191 352419
rect 126913 343449 127191 343727
rect 126913 325449 127191 325727
rect 126913 307449 127191 307727
rect 126913 289449 127191 289727
rect 126913 271449 127191 271727
rect 126913 253449 127191 253727
rect 126913 235449 127191 235727
rect 126913 217449 127191 217727
rect 126913 199449 127191 199727
rect 126913 181449 127191 181727
rect 126913 163449 127191 163727
rect 126913 145449 127191 145727
rect 126913 127449 127191 127727
rect 126913 109449 127191 109727
rect 126913 91449 127191 91727
rect 126913 73449 127191 73727
rect 126913 55449 127191 55727
rect 126913 37449 127191 37727
rect 126913 19449 127191 19727
rect 126913 1449 127191 1727
rect 126913 -451 127191 -173
rect 128773 345309 129051 345587
rect 128773 327309 129051 327587
rect 128773 309309 129051 309587
rect 128773 291309 129051 291587
rect 128773 273309 129051 273587
rect 128773 255309 129051 255587
rect 128773 237309 129051 237587
rect 128773 219309 129051 219587
rect 128773 201309 129051 201587
rect 128773 183309 129051 183587
rect 128773 165309 129051 165587
rect 128773 147309 129051 147587
rect 128773 129309 129051 129587
rect 128773 111309 129051 111587
rect 128773 93309 129051 93587
rect 128773 75309 129051 75587
rect 128773 57309 129051 57587
rect 128773 39309 129051 39587
rect 128773 21309 129051 21587
rect 128773 3309 129051 3587
rect 128773 -1411 129051 -1133
rect 130633 347169 130911 347447
rect 130633 329169 130911 329447
rect 130633 311169 130911 311447
rect 130633 293169 130911 293447
rect 130633 275169 130911 275447
rect 130633 257169 130911 257447
rect 130633 239169 130911 239447
rect 130633 221169 130911 221447
rect 130633 203169 130911 203447
rect 130633 185169 130911 185447
rect 130633 167169 130911 167447
rect 130633 149169 130911 149447
rect 130633 131169 130911 131447
rect 130633 113169 130911 113447
rect 130633 95169 130911 95447
rect 130633 77169 130911 77447
rect 130633 59169 130911 59447
rect 130633 41169 130911 41447
rect 130633 23169 130911 23447
rect 130633 5169 130911 5447
rect 130633 -2371 130911 -2093
rect 141493 355501 141771 355779
rect 139633 354541 139911 354819
rect 137773 353581 138051 353859
rect 132493 349029 132771 349307
rect 132493 331029 132771 331307
rect 132493 313029 132771 313307
rect 132493 295029 132771 295307
rect 132493 277029 132771 277307
rect 132493 259029 132771 259307
rect 132493 241029 132771 241307
rect 132493 223029 132771 223307
rect 132493 205029 132771 205307
rect 132493 187029 132771 187307
rect 132493 169029 132771 169307
rect 132493 151029 132771 151307
rect 132493 133029 132771 133307
rect 132493 115029 132771 115307
rect 132493 97029 132771 97307
rect 132493 79029 132771 79307
rect 132493 61029 132771 61307
rect 132493 43029 132771 43307
rect 132493 25029 132771 25307
rect 132493 7029 132771 7307
rect 123493 -3811 123771 -3533
rect 135913 352621 136191 352899
rect 135913 334449 136191 334727
rect 135913 316449 136191 316727
rect 135913 298449 136191 298727
rect 135913 280449 136191 280727
rect 135913 262449 136191 262727
rect 135913 244449 136191 244727
rect 135913 226449 136191 226727
rect 135913 208449 136191 208727
rect 135913 190449 136191 190727
rect 135913 172449 136191 172727
rect 135913 154449 136191 154727
rect 135913 136449 136191 136727
rect 135913 118449 136191 118727
rect 135913 100449 136191 100727
rect 135913 82449 136191 82727
rect 135913 64449 136191 64727
rect 135913 46449 136191 46727
rect 135913 28449 136191 28727
rect 135913 10449 136191 10727
rect 135913 -931 136191 -653
rect 137773 336309 138051 336587
rect 137773 318309 138051 318587
rect 137773 300309 138051 300587
rect 137773 282309 138051 282587
rect 137773 264309 138051 264587
rect 137773 246309 138051 246587
rect 137773 228309 138051 228587
rect 137773 210309 138051 210587
rect 137773 192309 138051 192587
rect 137773 174309 138051 174587
rect 137773 156309 138051 156587
rect 137773 138309 138051 138587
rect 137773 120309 138051 120587
rect 137773 102309 138051 102587
rect 137773 84309 138051 84587
rect 137773 66309 138051 66587
rect 137773 48309 138051 48587
rect 137773 30309 138051 30587
rect 137773 12309 138051 12587
rect 137773 -1891 138051 -1613
rect 139633 338169 139911 338447
rect 139633 320169 139911 320447
rect 139633 302169 139911 302447
rect 139633 284169 139911 284447
rect 139633 266169 139911 266447
rect 139633 248169 139911 248447
rect 139633 230169 139911 230447
rect 139633 212169 139911 212447
rect 139633 194169 139911 194447
rect 139633 176169 139911 176447
rect 139633 158169 139911 158447
rect 139633 140169 139911 140447
rect 139633 122169 139911 122447
rect 139633 104169 139911 104447
rect 139633 86169 139911 86447
rect 139633 68169 139911 68447
rect 139633 50169 139911 50447
rect 139633 32169 139911 32447
rect 139633 14169 139911 14447
rect 139633 -2851 139911 -2573
rect 150493 355021 150771 355299
rect 148633 354061 148911 354339
rect 146773 353101 147051 353379
rect 141493 340029 141771 340307
rect 141493 322029 141771 322307
rect 141493 304029 141771 304307
rect 141493 286029 141771 286307
rect 141493 268029 141771 268307
rect 141493 250029 141771 250307
rect 141493 232029 141771 232307
rect 141493 214029 141771 214307
rect 141493 196029 141771 196307
rect 141493 178029 141771 178307
rect 141493 160029 141771 160307
rect 141493 142029 141771 142307
rect 141493 124029 141771 124307
rect 141493 106029 141771 106307
rect 141493 88029 141771 88307
rect 141493 70029 141771 70307
rect 141493 52029 141771 52307
rect 141493 34029 141771 34307
rect 141493 16029 141771 16307
rect 132493 -3331 132771 -3053
rect 144913 352141 145191 352419
rect 144913 343449 145191 343727
rect 144913 325449 145191 325727
rect 144913 307449 145191 307727
rect 144913 289449 145191 289727
rect 144913 271449 145191 271727
rect 144913 253449 145191 253727
rect 144913 235449 145191 235727
rect 144913 217449 145191 217727
rect 144913 199449 145191 199727
rect 144913 181449 145191 181727
rect 144913 163449 145191 163727
rect 144913 145449 145191 145727
rect 144913 127449 145191 127727
rect 144913 109449 145191 109727
rect 144913 91449 145191 91727
rect 144913 73449 145191 73727
rect 144913 55449 145191 55727
rect 144913 37449 145191 37727
rect 144913 19449 145191 19727
rect 144913 1449 145191 1727
rect 144913 -451 145191 -173
rect 146773 345309 147051 345587
rect 146773 327309 147051 327587
rect 146773 309309 147051 309587
rect 146773 291309 147051 291587
rect 146773 273309 147051 273587
rect 146773 255309 147051 255587
rect 146773 237309 147051 237587
rect 146773 219309 147051 219587
rect 146773 201309 147051 201587
rect 146773 183309 147051 183587
rect 146773 165309 147051 165587
rect 146773 147309 147051 147587
rect 146773 129309 147051 129587
rect 146773 111309 147051 111587
rect 146773 93309 147051 93587
rect 146773 75309 147051 75587
rect 146773 57309 147051 57587
rect 146773 39309 147051 39587
rect 146773 21309 147051 21587
rect 146773 3309 147051 3587
rect 146773 -1411 147051 -1133
rect 148633 347169 148911 347447
rect 148633 329169 148911 329447
rect 148633 311169 148911 311447
rect 148633 293169 148911 293447
rect 148633 275169 148911 275447
rect 148633 257169 148911 257447
rect 148633 239169 148911 239447
rect 148633 221169 148911 221447
rect 148633 203169 148911 203447
rect 148633 185169 148911 185447
rect 148633 167169 148911 167447
rect 148633 149169 148911 149447
rect 148633 131169 148911 131447
rect 148633 113169 148911 113447
rect 148633 95169 148911 95447
rect 148633 77169 148911 77447
rect 148633 59169 148911 59447
rect 148633 41169 148911 41447
rect 148633 23169 148911 23447
rect 148633 5169 148911 5447
rect 148633 -2371 148911 -2093
rect 159493 355501 159771 355779
rect 157633 354541 157911 354819
rect 155773 353581 156051 353859
rect 150493 349029 150771 349307
rect 150493 331029 150771 331307
rect 150493 313029 150771 313307
rect 150493 295029 150771 295307
rect 150493 277029 150771 277307
rect 150493 259029 150771 259307
rect 150493 241029 150771 241307
rect 150493 223029 150771 223307
rect 150493 205029 150771 205307
rect 150493 187029 150771 187307
rect 150493 169029 150771 169307
rect 150493 151029 150771 151307
rect 150493 133029 150771 133307
rect 150493 115029 150771 115307
rect 150493 97029 150771 97307
rect 150493 79029 150771 79307
rect 150493 61029 150771 61307
rect 150493 43029 150771 43307
rect 150493 25029 150771 25307
rect 150493 7029 150771 7307
rect 141493 -3811 141771 -3533
rect 153913 352621 154191 352899
rect 153913 334449 154191 334727
rect 153913 316449 154191 316727
rect 153913 298449 154191 298727
rect 153913 280449 154191 280727
rect 153913 262449 154191 262727
rect 153913 244449 154191 244727
rect 153913 226449 154191 226727
rect 153913 208449 154191 208727
rect 153913 190449 154191 190727
rect 153913 172449 154191 172727
rect 153913 154449 154191 154727
rect 153913 136449 154191 136727
rect 153913 118449 154191 118727
rect 153913 100449 154191 100727
rect 153913 82449 154191 82727
rect 153913 64449 154191 64727
rect 153913 46449 154191 46727
rect 153913 28449 154191 28727
rect 153913 10449 154191 10727
rect 153913 -931 154191 -653
rect 155773 336309 156051 336587
rect 155773 318309 156051 318587
rect 155773 300309 156051 300587
rect 155773 282309 156051 282587
rect 155773 264309 156051 264587
rect 155773 246309 156051 246587
rect 155773 228309 156051 228587
rect 155773 210309 156051 210587
rect 155773 192309 156051 192587
rect 155773 174309 156051 174587
rect 155773 156309 156051 156587
rect 155773 138309 156051 138587
rect 155773 120309 156051 120587
rect 155773 102309 156051 102587
rect 155773 84309 156051 84587
rect 155773 66309 156051 66587
rect 155773 48309 156051 48587
rect 155773 30309 156051 30587
rect 155773 12309 156051 12587
rect 155773 -1891 156051 -1613
rect 157633 338169 157911 338447
rect 157633 320169 157911 320447
rect 157633 302169 157911 302447
rect 157633 284169 157911 284447
rect 157633 266169 157911 266447
rect 157633 248169 157911 248447
rect 157633 230169 157911 230447
rect 157633 212169 157911 212447
rect 157633 194169 157911 194447
rect 157633 176169 157911 176447
rect 157633 158169 157911 158447
rect 157633 140169 157911 140447
rect 157633 122169 157911 122447
rect 157633 104169 157911 104447
rect 157633 86169 157911 86447
rect 157633 68169 157911 68447
rect 157633 50169 157911 50447
rect 157633 32169 157911 32447
rect 157633 14169 157911 14447
rect 157633 -2851 157911 -2573
rect 168493 355021 168771 355299
rect 166633 354061 166911 354339
rect 164773 353101 165051 353379
rect 159493 340029 159771 340307
rect 159493 322029 159771 322307
rect 159493 304029 159771 304307
rect 159493 286029 159771 286307
rect 159493 268029 159771 268307
rect 159493 250029 159771 250307
rect 159493 232029 159771 232307
rect 159493 214029 159771 214307
rect 159493 196029 159771 196307
rect 159493 178029 159771 178307
rect 159493 160029 159771 160307
rect 159493 142029 159771 142307
rect 159493 124029 159771 124307
rect 159493 106029 159771 106307
rect 159493 88029 159771 88307
rect 159493 70029 159771 70307
rect 159493 52029 159771 52307
rect 159493 34029 159771 34307
rect 159493 16029 159771 16307
rect 150493 -3331 150771 -3053
rect 162913 352141 163191 352419
rect 162913 343449 163191 343727
rect 162913 325449 163191 325727
rect 162913 307449 163191 307727
rect 162913 289449 163191 289727
rect 162913 271449 163191 271727
rect 162913 253449 163191 253727
rect 162913 235449 163191 235727
rect 162913 217449 163191 217727
rect 162913 199449 163191 199727
rect 162913 181449 163191 181727
rect 162913 163449 163191 163727
rect 162913 145449 163191 145727
rect 162913 127449 163191 127727
rect 162913 109449 163191 109727
rect 162913 91449 163191 91727
rect 162913 73449 163191 73727
rect 162913 55449 163191 55727
rect 162913 37449 163191 37727
rect 162913 19449 163191 19727
rect 162913 1449 163191 1727
rect 162913 -451 163191 -173
rect 164773 345309 165051 345587
rect 164773 327309 165051 327587
rect 164773 309309 165051 309587
rect 164773 291309 165051 291587
rect 164773 273309 165051 273587
rect 164773 255309 165051 255587
rect 164773 237309 165051 237587
rect 164773 219309 165051 219587
rect 164773 201309 165051 201587
rect 164773 183309 165051 183587
rect 164773 165309 165051 165587
rect 164773 147309 165051 147587
rect 164773 129309 165051 129587
rect 164773 111309 165051 111587
rect 164773 93309 165051 93587
rect 164773 75309 165051 75587
rect 164773 57309 165051 57587
rect 164773 39309 165051 39587
rect 164773 21309 165051 21587
rect 164773 3309 165051 3587
rect 164773 -1411 165051 -1133
rect 166633 347169 166911 347447
rect 166633 329169 166911 329447
rect 166633 311169 166911 311447
rect 166633 293169 166911 293447
rect 166633 275169 166911 275447
rect 166633 257169 166911 257447
rect 166633 239169 166911 239447
rect 166633 221169 166911 221447
rect 166633 203169 166911 203447
rect 166633 185169 166911 185447
rect 166633 167169 166911 167447
rect 166633 149169 166911 149447
rect 166633 131169 166911 131447
rect 166633 113169 166911 113447
rect 166633 95169 166911 95447
rect 166633 77169 166911 77447
rect 166633 59169 166911 59447
rect 166633 41169 166911 41447
rect 166633 23169 166911 23447
rect 166633 5169 166911 5447
rect 166633 -2371 166911 -2093
rect 177493 355501 177771 355779
rect 175633 354541 175911 354819
rect 173773 353581 174051 353859
rect 168493 349029 168771 349307
rect 168493 331029 168771 331307
rect 168493 313029 168771 313307
rect 168493 295029 168771 295307
rect 168493 277029 168771 277307
rect 168493 259029 168771 259307
rect 168493 241029 168771 241307
rect 168493 223029 168771 223307
rect 168493 205029 168771 205307
rect 168493 187029 168771 187307
rect 168493 169029 168771 169307
rect 168493 151029 168771 151307
rect 168493 133029 168771 133307
rect 168493 115029 168771 115307
rect 168493 97029 168771 97307
rect 168493 79029 168771 79307
rect 168493 61029 168771 61307
rect 168493 43029 168771 43307
rect 168493 25029 168771 25307
rect 168493 7029 168771 7307
rect 159493 -3811 159771 -3533
rect 171913 352621 172191 352899
rect 171913 334449 172191 334727
rect 171913 316449 172191 316727
rect 171913 298449 172191 298727
rect 171913 280449 172191 280727
rect 171913 262449 172191 262727
rect 171913 244449 172191 244727
rect 171913 226449 172191 226727
rect 171913 208449 172191 208727
rect 171913 190449 172191 190727
rect 171913 172449 172191 172727
rect 171913 154449 172191 154727
rect 171913 136449 172191 136727
rect 171913 118449 172191 118727
rect 171913 100449 172191 100727
rect 171913 82449 172191 82727
rect 171913 64449 172191 64727
rect 171913 46449 172191 46727
rect 171913 28449 172191 28727
rect 171913 10449 172191 10727
rect 171913 -931 172191 -653
rect 173773 336309 174051 336587
rect 173773 318309 174051 318587
rect 173773 300309 174051 300587
rect 173773 282309 174051 282587
rect 173773 264309 174051 264587
rect 173773 246309 174051 246587
rect 173773 228309 174051 228587
rect 173773 210309 174051 210587
rect 173773 192309 174051 192587
rect 173773 174309 174051 174587
rect 173773 156309 174051 156587
rect 173773 138309 174051 138587
rect 173773 120309 174051 120587
rect 173773 102309 174051 102587
rect 173773 84309 174051 84587
rect 173773 66309 174051 66587
rect 173773 48309 174051 48587
rect 173773 30309 174051 30587
rect 173773 12309 174051 12587
rect 173773 -1891 174051 -1613
rect 175633 338169 175911 338447
rect 175633 320169 175911 320447
rect 175633 302169 175911 302447
rect 175633 284169 175911 284447
rect 175633 266169 175911 266447
rect 175633 248169 175911 248447
rect 175633 230169 175911 230447
rect 175633 212169 175911 212447
rect 175633 194169 175911 194447
rect 175633 176169 175911 176447
rect 175633 158169 175911 158447
rect 175633 140169 175911 140447
rect 175633 122169 175911 122447
rect 175633 104169 175911 104447
rect 175633 86169 175911 86447
rect 175633 68169 175911 68447
rect 175633 50169 175911 50447
rect 175633 32169 175911 32447
rect 175633 14169 175911 14447
rect 175633 -2851 175911 -2573
rect 186493 355021 186771 355299
rect 184633 354061 184911 354339
rect 182773 353101 183051 353379
rect 177493 340029 177771 340307
rect 177493 322029 177771 322307
rect 177493 304029 177771 304307
rect 177493 286029 177771 286307
rect 177493 268029 177771 268307
rect 177493 250029 177771 250307
rect 177493 232029 177771 232307
rect 177493 214029 177771 214307
rect 177493 196029 177771 196307
rect 177493 178029 177771 178307
rect 177493 160029 177771 160307
rect 177493 142029 177771 142307
rect 177493 124029 177771 124307
rect 177493 106029 177771 106307
rect 177493 88029 177771 88307
rect 177493 70029 177771 70307
rect 177493 52029 177771 52307
rect 177493 34029 177771 34307
rect 177493 16029 177771 16307
rect 168493 -3331 168771 -3053
rect 180913 352141 181191 352419
rect 180913 343449 181191 343727
rect 180913 325449 181191 325727
rect 180913 307449 181191 307727
rect 180913 289449 181191 289727
rect 180913 271449 181191 271727
rect 180913 253449 181191 253727
rect 180913 235449 181191 235727
rect 180913 217449 181191 217727
rect 180913 199449 181191 199727
rect 180913 181449 181191 181727
rect 180913 163449 181191 163727
rect 180913 145449 181191 145727
rect 180913 127449 181191 127727
rect 180913 109449 181191 109727
rect 180913 91449 181191 91727
rect 180913 73449 181191 73727
rect 180913 55449 181191 55727
rect 180913 37449 181191 37727
rect 180913 19449 181191 19727
rect 180913 1449 181191 1727
rect 180913 -451 181191 -173
rect 182773 345309 183051 345587
rect 182773 327309 183051 327587
rect 182773 309309 183051 309587
rect 182773 291309 183051 291587
rect 182773 273309 183051 273587
rect 182773 255309 183051 255587
rect 182773 237309 183051 237587
rect 182773 219309 183051 219587
rect 182773 201309 183051 201587
rect 182773 183309 183051 183587
rect 182773 165309 183051 165587
rect 182773 147309 183051 147587
rect 182773 129309 183051 129587
rect 182773 111309 183051 111587
rect 182773 93309 183051 93587
rect 182773 75309 183051 75587
rect 182773 57309 183051 57587
rect 182773 39309 183051 39587
rect 182773 21309 183051 21587
rect 182773 3309 183051 3587
rect 182773 -1411 183051 -1133
rect 184633 347169 184911 347447
rect 184633 329169 184911 329447
rect 184633 311169 184911 311447
rect 184633 293169 184911 293447
rect 184633 275169 184911 275447
rect 184633 257169 184911 257447
rect 184633 239169 184911 239447
rect 184633 221169 184911 221447
rect 184633 203169 184911 203447
rect 184633 185169 184911 185447
rect 184633 167169 184911 167447
rect 184633 149169 184911 149447
rect 184633 131169 184911 131447
rect 184633 113169 184911 113447
rect 184633 95169 184911 95447
rect 184633 77169 184911 77447
rect 184633 59169 184911 59447
rect 184633 41169 184911 41447
rect 184633 23169 184911 23447
rect 184633 5169 184911 5447
rect 184633 -2371 184911 -2093
rect 195493 355501 195771 355779
rect 193633 354541 193911 354819
rect 191773 353581 192051 353859
rect 186493 349029 186771 349307
rect 186493 331029 186771 331307
rect 186493 313029 186771 313307
rect 186493 295029 186771 295307
rect 186493 277029 186771 277307
rect 186493 259029 186771 259307
rect 186493 241029 186771 241307
rect 186493 223029 186771 223307
rect 186493 205029 186771 205307
rect 186493 187029 186771 187307
rect 186493 169029 186771 169307
rect 186493 151029 186771 151307
rect 186493 133029 186771 133307
rect 186493 115029 186771 115307
rect 186493 97029 186771 97307
rect 186493 79029 186771 79307
rect 186493 61029 186771 61307
rect 186493 43029 186771 43307
rect 186493 25029 186771 25307
rect 186493 7029 186771 7307
rect 177493 -3811 177771 -3533
rect 189913 352621 190191 352899
rect 189913 334449 190191 334727
rect 189913 316449 190191 316727
rect 189913 298449 190191 298727
rect 189913 280449 190191 280727
rect 189913 262449 190191 262727
rect 189913 244449 190191 244727
rect 189913 226449 190191 226727
rect 189913 208449 190191 208727
rect 189913 190449 190191 190727
rect 189913 172449 190191 172727
rect 189913 154449 190191 154727
rect 189913 136449 190191 136727
rect 189913 118449 190191 118727
rect 189913 100449 190191 100727
rect 189913 82449 190191 82727
rect 189913 64449 190191 64727
rect 189913 46449 190191 46727
rect 189913 28449 190191 28727
rect 189913 10449 190191 10727
rect 189913 -931 190191 -653
rect 191773 336309 192051 336587
rect 191773 318309 192051 318587
rect 191773 300309 192051 300587
rect 191773 282309 192051 282587
rect 191773 264309 192051 264587
rect 191773 246309 192051 246587
rect 191773 228309 192051 228587
rect 191773 210309 192051 210587
rect 191773 192309 192051 192587
rect 191773 174309 192051 174587
rect 191773 156309 192051 156587
rect 191773 138309 192051 138587
rect 191773 120309 192051 120587
rect 191773 102309 192051 102587
rect 191773 84309 192051 84587
rect 191773 66309 192051 66587
rect 191773 48309 192051 48587
rect 191773 30309 192051 30587
rect 191773 12309 192051 12587
rect 191773 -1891 192051 -1613
rect 193633 338169 193911 338447
rect 193633 320169 193911 320447
rect 193633 302169 193911 302447
rect 193633 284169 193911 284447
rect 193633 266169 193911 266447
rect 193633 248169 193911 248447
rect 193633 230169 193911 230447
rect 193633 212169 193911 212447
rect 193633 194169 193911 194447
rect 193633 176169 193911 176447
rect 193633 158169 193911 158447
rect 193633 140169 193911 140447
rect 193633 122169 193911 122447
rect 193633 104169 193911 104447
rect 193633 86169 193911 86447
rect 193633 68169 193911 68447
rect 193633 50169 193911 50447
rect 193633 32169 193911 32447
rect 193633 14169 193911 14447
rect 193633 -2851 193911 -2573
rect 204493 355021 204771 355299
rect 202633 354061 202911 354339
rect 200773 353101 201051 353379
rect 195493 340029 195771 340307
rect 195493 322029 195771 322307
rect 195493 304029 195771 304307
rect 195493 286029 195771 286307
rect 195493 268029 195771 268307
rect 195493 250029 195771 250307
rect 195493 232029 195771 232307
rect 195493 214029 195771 214307
rect 195493 196029 195771 196307
rect 195493 178029 195771 178307
rect 195493 160029 195771 160307
rect 195493 142029 195771 142307
rect 195493 124029 195771 124307
rect 195493 106029 195771 106307
rect 195493 88029 195771 88307
rect 195493 70029 195771 70307
rect 195493 52029 195771 52307
rect 195493 34029 195771 34307
rect 195493 16029 195771 16307
rect 186493 -3331 186771 -3053
rect 198913 352141 199191 352419
rect 198913 343449 199191 343727
rect 198913 325449 199191 325727
rect 198913 307449 199191 307727
rect 198913 289449 199191 289727
rect 198913 271449 199191 271727
rect 198913 253449 199191 253727
rect 198913 235449 199191 235727
rect 198913 217449 199191 217727
rect 198913 199449 199191 199727
rect 198913 181449 199191 181727
rect 198913 163449 199191 163727
rect 198913 145449 199191 145727
rect 198913 127449 199191 127727
rect 198913 109449 199191 109727
rect 198913 91449 199191 91727
rect 198913 73449 199191 73727
rect 198913 55449 199191 55727
rect 198913 37449 199191 37727
rect 198913 19449 199191 19727
rect 198913 1449 199191 1727
rect 198913 -451 199191 -173
rect 200773 345309 201051 345587
rect 200773 327309 201051 327587
rect 200773 309309 201051 309587
rect 200773 291309 201051 291587
rect 200773 273309 201051 273587
rect 200773 255309 201051 255587
rect 200773 237309 201051 237587
rect 200773 219309 201051 219587
rect 200773 201309 201051 201587
rect 200773 183309 201051 183587
rect 200773 165309 201051 165587
rect 200773 147309 201051 147587
rect 200773 129309 201051 129587
rect 200773 111309 201051 111587
rect 200773 93309 201051 93587
rect 200773 75309 201051 75587
rect 200773 57309 201051 57587
rect 200773 39309 201051 39587
rect 200773 21309 201051 21587
rect 200773 3309 201051 3587
rect 200773 -1411 201051 -1133
rect 202633 347169 202911 347447
rect 202633 329169 202911 329447
rect 202633 311169 202911 311447
rect 202633 293169 202911 293447
rect 202633 275169 202911 275447
rect 202633 257169 202911 257447
rect 202633 239169 202911 239447
rect 202633 221169 202911 221447
rect 202633 203169 202911 203447
rect 202633 185169 202911 185447
rect 202633 167169 202911 167447
rect 202633 149169 202911 149447
rect 202633 131169 202911 131447
rect 202633 113169 202911 113447
rect 202633 95169 202911 95447
rect 202633 77169 202911 77447
rect 202633 59169 202911 59447
rect 202633 41169 202911 41447
rect 202633 23169 202911 23447
rect 202633 5169 202911 5447
rect 202633 -2371 202911 -2093
rect 213493 355501 213771 355779
rect 211633 354541 211911 354819
rect 209773 353581 210051 353859
rect 204493 349029 204771 349307
rect 204493 331029 204771 331307
rect 204493 313029 204771 313307
rect 204493 295029 204771 295307
rect 204493 277029 204771 277307
rect 204493 259029 204771 259307
rect 204493 241029 204771 241307
rect 204493 223029 204771 223307
rect 204493 205029 204771 205307
rect 204493 187029 204771 187307
rect 204493 169029 204771 169307
rect 204493 151029 204771 151307
rect 204493 133029 204771 133307
rect 204493 115029 204771 115307
rect 204493 97029 204771 97307
rect 204493 79029 204771 79307
rect 204493 61029 204771 61307
rect 204493 43029 204771 43307
rect 204493 25029 204771 25307
rect 204493 7029 204771 7307
rect 195493 -3811 195771 -3533
rect 207913 352621 208191 352899
rect 207913 334449 208191 334727
rect 207913 316449 208191 316727
rect 207913 298449 208191 298727
rect 207913 280449 208191 280727
rect 207913 262449 208191 262727
rect 207913 244449 208191 244727
rect 207913 226449 208191 226727
rect 207913 208449 208191 208727
rect 207913 190449 208191 190727
rect 207913 172449 208191 172727
rect 207913 154449 208191 154727
rect 207913 136449 208191 136727
rect 207913 118449 208191 118727
rect 207913 100449 208191 100727
rect 207913 82449 208191 82727
rect 207913 64449 208191 64727
rect 207913 46449 208191 46727
rect 207913 28449 208191 28727
rect 207913 10449 208191 10727
rect 207913 -931 208191 -653
rect 209773 336309 210051 336587
rect 209773 318309 210051 318587
rect 209773 300309 210051 300587
rect 209773 282309 210051 282587
rect 209773 264309 210051 264587
rect 209773 246309 210051 246587
rect 209773 228309 210051 228587
rect 209773 210309 210051 210587
rect 209773 192309 210051 192587
rect 209773 174309 210051 174587
rect 209773 156309 210051 156587
rect 209773 138309 210051 138587
rect 209773 120309 210051 120587
rect 209773 102309 210051 102587
rect 209773 84309 210051 84587
rect 209773 66309 210051 66587
rect 209773 48309 210051 48587
rect 209773 30309 210051 30587
rect 209773 12309 210051 12587
rect 209773 -1891 210051 -1613
rect 211633 338169 211911 338447
rect 211633 320169 211911 320447
rect 211633 302169 211911 302447
rect 211633 284169 211911 284447
rect 211633 266169 211911 266447
rect 211633 248169 211911 248447
rect 211633 230169 211911 230447
rect 211633 212169 211911 212447
rect 211633 194169 211911 194447
rect 211633 176169 211911 176447
rect 211633 158169 211911 158447
rect 211633 140169 211911 140447
rect 211633 122169 211911 122447
rect 211633 104169 211911 104447
rect 211633 86169 211911 86447
rect 211633 68169 211911 68447
rect 211633 50169 211911 50447
rect 211633 32169 211911 32447
rect 211633 14169 211911 14447
rect 211633 -2851 211911 -2573
rect 222493 355021 222771 355299
rect 220633 354061 220911 354339
rect 218773 353101 219051 353379
rect 213493 340029 213771 340307
rect 213493 322029 213771 322307
rect 213493 304029 213771 304307
rect 213493 286029 213771 286307
rect 213493 268029 213771 268307
rect 213493 250029 213771 250307
rect 213493 232029 213771 232307
rect 213493 214029 213771 214307
rect 213493 196029 213771 196307
rect 213493 178029 213771 178307
rect 213493 160029 213771 160307
rect 213493 142029 213771 142307
rect 213493 124029 213771 124307
rect 213493 106029 213771 106307
rect 213493 88029 213771 88307
rect 213493 70029 213771 70307
rect 213493 52029 213771 52307
rect 213493 34029 213771 34307
rect 213493 16029 213771 16307
rect 204493 -3331 204771 -3053
rect 216913 352141 217191 352419
rect 216913 343449 217191 343727
rect 216913 325449 217191 325727
rect 216913 307449 217191 307727
rect 216913 289449 217191 289727
rect 216913 271449 217191 271727
rect 216913 253449 217191 253727
rect 216913 235449 217191 235727
rect 216913 217449 217191 217727
rect 216913 199449 217191 199727
rect 216913 181449 217191 181727
rect 216913 163449 217191 163727
rect 216913 145449 217191 145727
rect 216913 127449 217191 127727
rect 216913 109449 217191 109727
rect 216913 91449 217191 91727
rect 216913 73449 217191 73727
rect 216913 55449 217191 55727
rect 216913 37449 217191 37727
rect 216913 19449 217191 19727
rect 216913 1449 217191 1727
rect 216913 -451 217191 -173
rect 218773 345309 219051 345587
rect 218773 327309 219051 327587
rect 218773 309309 219051 309587
rect 218773 291309 219051 291587
rect 218773 273309 219051 273587
rect 218773 255309 219051 255587
rect 218773 237309 219051 237587
rect 218773 219309 219051 219587
rect 218773 201309 219051 201587
rect 218773 183309 219051 183587
rect 218773 165309 219051 165587
rect 218773 147309 219051 147587
rect 218773 129309 219051 129587
rect 218773 111309 219051 111587
rect 218773 93309 219051 93587
rect 218773 75309 219051 75587
rect 218773 57309 219051 57587
rect 218773 39309 219051 39587
rect 218773 21309 219051 21587
rect 218773 3309 219051 3587
rect 218773 -1411 219051 -1133
rect 220633 347169 220911 347447
rect 220633 329169 220911 329447
rect 220633 311169 220911 311447
rect 220633 293169 220911 293447
rect 220633 275169 220911 275447
rect 220633 257169 220911 257447
rect 220633 239169 220911 239447
rect 220633 221169 220911 221447
rect 220633 203169 220911 203447
rect 220633 185169 220911 185447
rect 220633 167169 220911 167447
rect 220633 149169 220911 149447
rect 220633 131169 220911 131447
rect 220633 113169 220911 113447
rect 220633 95169 220911 95447
rect 220633 77169 220911 77447
rect 220633 59169 220911 59447
rect 220633 41169 220911 41447
rect 220633 23169 220911 23447
rect 220633 5169 220911 5447
rect 220633 -2371 220911 -2093
rect 231493 355501 231771 355779
rect 229633 354541 229911 354819
rect 227773 353581 228051 353859
rect 222493 349029 222771 349307
rect 222493 331029 222771 331307
rect 222493 313029 222771 313307
rect 222493 295029 222771 295307
rect 222493 277029 222771 277307
rect 222493 259029 222771 259307
rect 222493 241029 222771 241307
rect 222493 223029 222771 223307
rect 222493 205029 222771 205307
rect 222493 187029 222771 187307
rect 222493 169029 222771 169307
rect 222493 151029 222771 151307
rect 222493 133029 222771 133307
rect 222493 115029 222771 115307
rect 222493 97029 222771 97307
rect 222493 79029 222771 79307
rect 222493 61029 222771 61307
rect 222493 43029 222771 43307
rect 222493 25029 222771 25307
rect 222493 7029 222771 7307
rect 213493 -3811 213771 -3533
rect 225913 352621 226191 352899
rect 225913 334449 226191 334727
rect 225913 316449 226191 316727
rect 225913 298449 226191 298727
rect 225913 280449 226191 280727
rect 225913 262449 226191 262727
rect 225913 244449 226191 244727
rect 225913 226449 226191 226727
rect 225913 208449 226191 208727
rect 225913 190449 226191 190727
rect 225913 172449 226191 172727
rect 225913 154449 226191 154727
rect 225913 136449 226191 136727
rect 225913 118449 226191 118727
rect 225913 100449 226191 100727
rect 225913 82449 226191 82727
rect 225913 64449 226191 64727
rect 225913 46449 226191 46727
rect 225913 28449 226191 28727
rect 225913 10449 226191 10727
rect 225913 -931 226191 -653
rect 227773 336309 228051 336587
rect 227773 318309 228051 318587
rect 227773 300309 228051 300587
rect 227773 282309 228051 282587
rect 227773 264309 228051 264587
rect 227773 246309 228051 246587
rect 227773 228309 228051 228587
rect 227773 210309 228051 210587
rect 227773 192309 228051 192587
rect 227773 174309 228051 174587
rect 227773 156309 228051 156587
rect 227773 138309 228051 138587
rect 227773 120309 228051 120587
rect 227773 102309 228051 102587
rect 227773 84309 228051 84587
rect 227773 66309 228051 66587
rect 227773 48309 228051 48587
rect 227773 30309 228051 30587
rect 227773 12309 228051 12587
rect 227773 -1891 228051 -1613
rect 229633 338169 229911 338447
rect 229633 320169 229911 320447
rect 229633 302169 229911 302447
rect 229633 284169 229911 284447
rect 229633 266169 229911 266447
rect 229633 248169 229911 248447
rect 229633 230169 229911 230447
rect 229633 212169 229911 212447
rect 229633 194169 229911 194447
rect 229633 176169 229911 176447
rect 229633 158169 229911 158447
rect 229633 140169 229911 140447
rect 229633 122169 229911 122447
rect 229633 104169 229911 104447
rect 229633 86169 229911 86447
rect 229633 68169 229911 68447
rect 229633 50169 229911 50447
rect 229633 32169 229911 32447
rect 229633 14169 229911 14447
rect 229633 -2851 229911 -2573
rect 240493 355021 240771 355299
rect 238633 354061 238911 354339
rect 236773 353101 237051 353379
rect 231493 340029 231771 340307
rect 231493 322029 231771 322307
rect 231493 304029 231771 304307
rect 231493 286029 231771 286307
rect 231493 268029 231771 268307
rect 231493 250029 231771 250307
rect 231493 232029 231771 232307
rect 231493 214029 231771 214307
rect 231493 196029 231771 196307
rect 231493 178029 231771 178307
rect 231493 160029 231771 160307
rect 231493 142029 231771 142307
rect 231493 124029 231771 124307
rect 231493 106029 231771 106307
rect 231493 88029 231771 88307
rect 231493 70029 231771 70307
rect 231493 52029 231771 52307
rect 231493 34029 231771 34307
rect 231493 16029 231771 16307
rect 222493 -3331 222771 -3053
rect 234913 352141 235191 352419
rect 234913 343449 235191 343727
rect 234913 325449 235191 325727
rect 234913 307449 235191 307727
rect 234913 289449 235191 289727
rect 234913 271449 235191 271727
rect 234913 253449 235191 253727
rect 234913 235449 235191 235727
rect 234913 217449 235191 217727
rect 234913 199449 235191 199727
rect 234913 181449 235191 181727
rect 234913 163449 235191 163727
rect 234913 145449 235191 145727
rect 234913 127449 235191 127727
rect 234913 109449 235191 109727
rect 234913 91449 235191 91727
rect 234913 73449 235191 73727
rect 234913 55449 235191 55727
rect 234913 37449 235191 37727
rect 234913 19449 235191 19727
rect 234913 1449 235191 1727
rect 234913 -451 235191 -173
rect 236773 345309 237051 345587
rect 236773 327309 237051 327587
rect 236773 309309 237051 309587
rect 236773 291309 237051 291587
rect 236773 273309 237051 273587
rect 236773 255309 237051 255587
rect 236773 237309 237051 237587
rect 236773 219309 237051 219587
rect 236773 201309 237051 201587
rect 236773 183309 237051 183587
rect 236773 165309 237051 165587
rect 236773 147309 237051 147587
rect 236773 129309 237051 129587
rect 236773 111309 237051 111587
rect 236773 93309 237051 93587
rect 236773 75309 237051 75587
rect 236773 57309 237051 57587
rect 236773 39309 237051 39587
rect 236773 21309 237051 21587
rect 236773 3309 237051 3587
rect 236773 -1411 237051 -1133
rect 238633 347169 238911 347447
rect 238633 329169 238911 329447
rect 238633 311169 238911 311447
rect 238633 293169 238911 293447
rect 238633 275169 238911 275447
rect 238633 257169 238911 257447
rect 238633 239169 238911 239447
rect 238633 221169 238911 221447
rect 238633 203169 238911 203447
rect 238633 185169 238911 185447
rect 238633 167169 238911 167447
rect 238633 149169 238911 149447
rect 238633 131169 238911 131447
rect 238633 113169 238911 113447
rect 238633 95169 238911 95447
rect 238633 77169 238911 77447
rect 238633 59169 238911 59447
rect 238633 41169 238911 41447
rect 238633 23169 238911 23447
rect 238633 5169 238911 5447
rect 238633 -2371 238911 -2093
rect 249493 355501 249771 355779
rect 247633 354541 247911 354819
rect 245773 353581 246051 353859
rect 240493 349029 240771 349307
rect 240493 331029 240771 331307
rect 240493 313029 240771 313307
rect 240493 295029 240771 295307
rect 240493 277029 240771 277307
rect 240493 259029 240771 259307
rect 240493 241029 240771 241307
rect 240493 223029 240771 223307
rect 240493 205029 240771 205307
rect 240493 187029 240771 187307
rect 240493 169029 240771 169307
rect 240493 151029 240771 151307
rect 240493 133029 240771 133307
rect 240493 115029 240771 115307
rect 240493 97029 240771 97307
rect 240493 79029 240771 79307
rect 240493 61029 240771 61307
rect 240493 43029 240771 43307
rect 240493 25029 240771 25307
rect 240493 7029 240771 7307
rect 231493 -3811 231771 -3533
rect 243913 352621 244191 352899
rect 243913 334449 244191 334727
rect 243913 316449 244191 316727
rect 243913 298449 244191 298727
rect 243913 280449 244191 280727
rect 243913 262449 244191 262727
rect 243913 244449 244191 244727
rect 243913 226449 244191 226727
rect 243913 208449 244191 208727
rect 243913 190449 244191 190727
rect 243913 172449 244191 172727
rect 243913 154449 244191 154727
rect 243913 136449 244191 136727
rect 243913 118449 244191 118727
rect 243913 100449 244191 100727
rect 243913 82449 244191 82727
rect 243913 64449 244191 64727
rect 243913 46449 244191 46727
rect 243913 28449 244191 28727
rect 243913 10449 244191 10727
rect 243913 -931 244191 -653
rect 245773 336309 246051 336587
rect 245773 318309 246051 318587
rect 245773 300309 246051 300587
rect 245773 282309 246051 282587
rect 245773 264309 246051 264587
rect 245773 246309 246051 246587
rect 245773 228309 246051 228587
rect 245773 210309 246051 210587
rect 245773 192309 246051 192587
rect 245773 174309 246051 174587
rect 245773 156309 246051 156587
rect 245773 138309 246051 138587
rect 245773 120309 246051 120587
rect 245773 102309 246051 102587
rect 245773 84309 246051 84587
rect 245773 66309 246051 66587
rect 245773 48309 246051 48587
rect 245773 30309 246051 30587
rect 245773 12309 246051 12587
rect 245773 -1891 246051 -1613
rect 247633 338169 247911 338447
rect 247633 320169 247911 320447
rect 247633 302169 247911 302447
rect 247633 284169 247911 284447
rect 247633 266169 247911 266447
rect 247633 248169 247911 248447
rect 247633 230169 247911 230447
rect 247633 212169 247911 212447
rect 247633 194169 247911 194447
rect 247633 176169 247911 176447
rect 247633 158169 247911 158447
rect 247633 140169 247911 140447
rect 247633 122169 247911 122447
rect 247633 104169 247911 104447
rect 247633 86169 247911 86447
rect 247633 68169 247911 68447
rect 247633 50169 247911 50447
rect 247633 32169 247911 32447
rect 247633 14169 247911 14447
rect 247633 -2851 247911 -2573
rect 258493 355021 258771 355299
rect 256633 354061 256911 354339
rect 254773 353101 255051 353379
rect 249493 340029 249771 340307
rect 249493 322029 249771 322307
rect 249493 304029 249771 304307
rect 249493 286029 249771 286307
rect 249493 268029 249771 268307
rect 249493 250029 249771 250307
rect 249493 232029 249771 232307
rect 249493 214029 249771 214307
rect 249493 196029 249771 196307
rect 249493 178029 249771 178307
rect 249493 160029 249771 160307
rect 249493 142029 249771 142307
rect 249493 124029 249771 124307
rect 249493 106029 249771 106307
rect 249493 88029 249771 88307
rect 249493 70029 249771 70307
rect 249493 52029 249771 52307
rect 249493 34029 249771 34307
rect 249493 16029 249771 16307
rect 240493 -3331 240771 -3053
rect 252913 352141 253191 352419
rect 252913 343449 253191 343727
rect 252913 325449 253191 325727
rect 252913 307449 253191 307727
rect 252913 289449 253191 289727
rect 252913 271449 253191 271727
rect 252913 253449 253191 253727
rect 252913 235449 253191 235727
rect 252913 217449 253191 217727
rect 252913 199449 253191 199727
rect 252913 181449 253191 181727
rect 252913 163449 253191 163727
rect 252913 145449 253191 145727
rect 252913 127449 253191 127727
rect 252913 109449 253191 109727
rect 252913 91449 253191 91727
rect 252913 73449 253191 73727
rect 252913 55449 253191 55727
rect 252913 37449 253191 37727
rect 252913 19449 253191 19727
rect 252913 1449 253191 1727
rect 252913 -451 253191 -173
rect 254773 345309 255051 345587
rect 254773 327309 255051 327587
rect 254773 309309 255051 309587
rect 254773 291309 255051 291587
rect 254773 273309 255051 273587
rect 254773 255309 255051 255587
rect 254773 237309 255051 237587
rect 254773 219309 255051 219587
rect 254773 201309 255051 201587
rect 254773 183309 255051 183587
rect 254773 165309 255051 165587
rect 254773 147309 255051 147587
rect 254773 129309 255051 129587
rect 254773 111309 255051 111587
rect 254773 93309 255051 93587
rect 254773 75309 255051 75587
rect 254773 57309 255051 57587
rect 254773 39309 255051 39587
rect 254773 21309 255051 21587
rect 254773 3309 255051 3587
rect 254773 -1411 255051 -1133
rect 256633 347169 256911 347447
rect 256633 329169 256911 329447
rect 256633 311169 256911 311447
rect 256633 293169 256911 293447
rect 256633 275169 256911 275447
rect 256633 257169 256911 257447
rect 256633 239169 256911 239447
rect 256633 221169 256911 221447
rect 256633 203169 256911 203447
rect 256633 185169 256911 185447
rect 256633 167169 256911 167447
rect 256633 149169 256911 149447
rect 256633 131169 256911 131447
rect 256633 113169 256911 113447
rect 256633 95169 256911 95447
rect 256633 77169 256911 77447
rect 256633 59169 256911 59447
rect 256633 41169 256911 41447
rect 256633 23169 256911 23447
rect 256633 5169 256911 5447
rect 256633 -2371 256911 -2093
rect 267493 355501 267771 355779
rect 265633 354541 265911 354819
rect 263773 353581 264051 353859
rect 258493 349029 258771 349307
rect 258493 331029 258771 331307
rect 258493 313029 258771 313307
rect 258493 295029 258771 295307
rect 258493 277029 258771 277307
rect 258493 259029 258771 259307
rect 258493 241029 258771 241307
rect 258493 223029 258771 223307
rect 258493 205029 258771 205307
rect 258493 187029 258771 187307
rect 258493 169029 258771 169307
rect 258493 151029 258771 151307
rect 258493 133029 258771 133307
rect 258493 115029 258771 115307
rect 258493 97029 258771 97307
rect 258493 79029 258771 79307
rect 258493 61029 258771 61307
rect 258493 43029 258771 43307
rect 258493 25029 258771 25307
rect 258493 7029 258771 7307
rect 249493 -3811 249771 -3533
rect 261913 352621 262191 352899
rect 261913 334449 262191 334727
rect 261913 316449 262191 316727
rect 261913 298449 262191 298727
rect 261913 280449 262191 280727
rect 261913 262449 262191 262727
rect 261913 244449 262191 244727
rect 261913 226449 262191 226727
rect 261913 208449 262191 208727
rect 261913 190449 262191 190727
rect 261913 172449 262191 172727
rect 261913 154449 262191 154727
rect 261913 136449 262191 136727
rect 261913 118449 262191 118727
rect 261913 100449 262191 100727
rect 261913 82449 262191 82727
rect 261913 64449 262191 64727
rect 261913 46449 262191 46727
rect 261913 28449 262191 28727
rect 261913 10449 262191 10727
rect 261913 -931 262191 -653
rect 263773 336309 264051 336587
rect 263773 318309 264051 318587
rect 263773 300309 264051 300587
rect 263773 282309 264051 282587
rect 263773 264309 264051 264587
rect 263773 246309 264051 246587
rect 263773 228309 264051 228587
rect 263773 210309 264051 210587
rect 263773 192309 264051 192587
rect 263773 174309 264051 174587
rect 263773 156309 264051 156587
rect 263773 138309 264051 138587
rect 263773 120309 264051 120587
rect 263773 102309 264051 102587
rect 263773 84309 264051 84587
rect 263773 66309 264051 66587
rect 263773 48309 264051 48587
rect 263773 30309 264051 30587
rect 263773 12309 264051 12587
rect 263773 -1891 264051 -1613
rect 265633 338169 265911 338447
rect 265633 320169 265911 320447
rect 265633 302169 265911 302447
rect 265633 284169 265911 284447
rect 265633 266169 265911 266447
rect 265633 248169 265911 248447
rect 265633 230169 265911 230447
rect 265633 212169 265911 212447
rect 265633 194169 265911 194447
rect 265633 176169 265911 176447
rect 265633 158169 265911 158447
rect 265633 140169 265911 140447
rect 265633 122169 265911 122447
rect 265633 104169 265911 104447
rect 265633 86169 265911 86447
rect 265633 68169 265911 68447
rect 265633 50169 265911 50447
rect 265633 32169 265911 32447
rect 265633 14169 265911 14447
rect 265633 -2851 265911 -2573
rect 276493 355021 276771 355299
rect 274633 354061 274911 354339
rect 272773 353101 273051 353379
rect 267493 340029 267771 340307
rect 267493 322029 267771 322307
rect 267493 304029 267771 304307
rect 267493 286029 267771 286307
rect 267493 268029 267771 268307
rect 267493 250029 267771 250307
rect 267493 232029 267771 232307
rect 267493 214029 267771 214307
rect 267493 196029 267771 196307
rect 267493 178029 267771 178307
rect 267493 160029 267771 160307
rect 267493 142029 267771 142307
rect 267493 124029 267771 124307
rect 267493 106029 267771 106307
rect 267493 88029 267771 88307
rect 267493 70029 267771 70307
rect 267493 52029 267771 52307
rect 267493 34029 267771 34307
rect 267493 16029 267771 16307
rect 258493 -3331 258771 -3053
rect 270913 352141 271191 352419
rect 270913 343449 271191 343727
rect 270913 325449 271191 325727
rect 270913 307449 271191 307727
rect 270913 289449 271191 289727
rect 270913 271449 271191 271727
rect 270913 253449 271191 253727
rect 270913 235449 271191 235727
rect 270913 217449 271191 217727
rect 270913 199449 271191 199727
rect 270913 181449 271191 181727
rect 270913 163449 271191 163727
rect 270913 145449 271191 145727
rect 270913 127449 271191 127727
rect 270913 109449 271191 109727
rect 270913 91449 271191 91727
rect 270913 73449 271191 73727
rect 270913 55449 271191 55727
rect 270913 37449 271191 37727
rect 270913 19449 271191 19727
rect 270913 1449 271191 1727
rect 270913 -451 271191 -173
rect 272773 345309 273051 345587
rect 272773 327309 273051 327587
rect 272773 309309 273051 309587
rect 272773 291309 273051 291587
rect 272773 273309 273051 273587
rect 272773 255309 273051 255587
rect 272773 237309 273051 237587
rect 272773 219309 273051 219587
rect 272773 201309 273051 201587
rect 272773 183309 273051 183587
rect 272773 165309 273051 165587
rect 272773 147309 273051 147587
rect 272773 129309 273051 129587
rect 272773 111309 273051 111587
rect 272773 93309 273051 93587
rect 272773 75309 273051 75587
rect 272773 57309 273051 57587
rect 272773 39309 273051 39587
rect 272773 21309 273051 21587
rect 272773 3309 273051 3587
rect 272773 -1411 273051 -1133
rect 274633 347169 274911 347447
rect 274633 329169 274911 329447
rect 274633 311169 274911 311447
rect 274633 293169 274911 293447
rect 274633 275169 274911 275447
rect 274633 257169 274911 257447
rect 274633 239169 274911 239447
rect 274633 221169 274911 221447
rect 274633 203169 274911 203447
rect 274633 185169 274911 185447
rect 274633 167169 274911 167447
rect 274633 149169 274911 149447
rect 274633 131169 274911 131447
rect 274633 113169 274911 113447
rect 274633 95169 274911 95447
rect 274633 77169 274911 77447
rect 274633 59169 274911 59447
rect 274633 41169 274911 41447
rect 274633 23169 274911 23447
rect 274633 5169 274911 5447
rect 274633 -2371 274911 -2093
rect 285493 355501 285771 355779
rect 283633 354541 283911 354819
rect 281773 353581 282051 353859
rect 276493 349029 276771 349307
rect 276493 331029 276771 331307
rect 276493 313029 276771 313307
rect 276493 295029 276771 295307
rect 276493 277029 276771 277307
rect 276493 259029 276771 259307
rect 276493 241029 276771 241307
rect 276493 223029 276771 223307
rect 276493 205029 276771 205307
rect 276493 187029 276771 187307
rect 276493 169029 276771 169307
rect 276493 151029 276771 151307
rect 276493 133029 276771 133307
rect 276493 115029 276771 115307
rect 276493 97029 276771 97307
rect 276493 79029 276771 79307
rect 276493 61029 276771 61307
rect 276493 43029 276771 43307
rect 276493 25029 276771 25307
rect 276493 7029 276771 7307
rect 267493 -3811 267771 -3533
rect 279913 352621 280191 352899
rect 279913 334449 280191 334727
rect 279913 316449 280191 316727
rect 279913 298449 280191 298727
rect 279913 280449 280191 280727
rect 279913 262449 280191 262727
rect 279913 244449 280191 244727
rect 279913 226449 280191 226727
rect 279913 208449 280191 208727
rect 279913 190449 280191 190727
rect 279913 172449 280191 172727
rect 279913 154449 280191 154727
rect 279913 136449 280191 136727
rect 279913 118449 280191 118727
rect 279913 100449 280191 100727
rect 279913 82449 280191 82727
rect 279913 64449 280191 64727
rect 279913 46449 280191 46727
rect 279913 28449 280191 28727
rect 279913 10449 280191 10727
rect 279913 -931 280191 -653
rect 281773 336309 282051 336587
rect 281773 318309 282051 318587
rect 281773 300309 282051 300587
rect 281773 282309 282051 282587
rect 281773 264309 282051 264587
rect 281773 246309 282051 246587
rect 281773 228309 282051 228587
rect 281773 210309 282051 210587
rect 281773 192309 282051 192587
rect 281773 174309 282051 174587
rect 281773 156309 282051 156587
rect 281773 138309 282051 138587
rect 281773 120309 282051 120587
rect 281773 102309 282051 102587
rect 281773 84309 282051 84587
rect 281773 66309 282051 66587
rect 281773 48309 282051 48587
rect 281773 30309 282051 30587
rect 281773 12309 282051 12587
rect 281773 -1891 282051 -1613
rect 283633 338169 283911 338447
rect 283633 320169 283911 320447
rect 283633 302169 283911 302447
rect 283633 284169 283911 284447
rect 283633 266169 283911 266447
rect 283633 248169 283911 248447
rect 283633 230169 283911 230447
rect 283633 212169 283911 212447
rect 283633 194169 283911 194447
rect 283633 176169 283911 176447
rect 283633 158169 283911 158447
rect 283633 140169 283911 140447
rect 283633 122169 283911 122447
rect 283633 104169 283911 104447
rect 283633 86169 283911 86447
rect 283633 68169 283911 68447
rect 283633 50169 283911 50447
rect 283633 32169 283911 32447
rect 283633 14169 283911 14447
rect 283633 -2851 283911 -2573
rect 296031 355501 296309 355779
rect 295551 355021 295829 355299
rect 295071 354541 295349 354819
rect 294591 354061 294869 354339
rect 294111 353581 294389 353859
rect 290773 353101 291051 353379
rect 285493 340029 285771 340307
rect 285493 322029 285771 322307
rect 285493 304029 285771 304307
rect 285493 286029 285771 286307
rect 285493 268029 285771 268307
rect 285493 250029 285771 250307
rect 285493 232029 285771 232307
rect 285493 214029 285771 214307
rect 285493 196029 285771 196307
rect 285493 178029 285771 178307
rect 285493 160029 285771 160307
rect 285493 142029 285771 142307
rect 285493 124029 285771 124307
rect 285493 106029 285771 106307
rect 285493 88029 285771 88307
rect 285493 70029 285771 70307
rect 285493 52029 285771 52307
rect 285493 34029 285771 34307
rect 285493 16029 285771 16307
rect 276493 -3331 276771 -3053
rect 288913 352141 289191 352419
rect 288913 343449 289191 343727
rect 288913 325449 289191 325727
rect 288913 307449 289191 307727
rect 288913 289449 289191 289727
rect 288913 271449 289191 271727
rect 288913 253449 289191 253727
rect 288913 235449 289191 235727
rect 288913 217449 289191 217727
rect 288913 199449 289191 199727
rect 288913 181449 289191 181727
rect 288913 163449 289191 163727
rect 288913 145449 289191 145727
rect 288913 127449 289191 127727
rect 288913 109449 289191 109727
rect 288913 91449 289191 91727
rect 288913 73449 289191 73727
rect 288913 55449 289191 55727
rect 288913 37449 289191 37727
rect 288913 19449 289191 19727
rect 288913 1449 289191 1727
rect 288913 -451 289191 -173
rect 293631 353101 293909 353379
rect 293151 352621 293429 352899
rect 290773 345309 291051 345587
rect 290773 327309 291051 327587
rect 290773 309309 291051 309587
rect 290773 291309 291051 291587
rect 290773 273309 291051 273587
rect 290773 255309 291051 255587
rect 290773 237309 291051 237587
rect 290773 219309 291051 219587
rect 290773 201309 291051 201587
rect 290773 183309 291051 183587
rect 290773 165309 291051 165587
rect 290773 147309 291051 147587
rect 290773 129309 291051 129587
rect 290773 111309 291051 111587
rect 290773 93309 291051 93587
rect 290773 75309 291051 75587
rect 290773 57309 291051 57587
rect 290773 39309 291051 39587
rect 290773 21309 291051 21587
rect 290773 3309 291051 3587
rect 292671 352141 292949 352419
rect 292671 343449 292949 343727
rect 292671 325449 292949 325727
rect 292671 307449 292949 307727
rect 292671 289449 292949 289727
rect 292671 271449 292949 271727
rect 292671 253449 292949 253727
rect 292671 235449 292949 235727
rect 292671 217449 292949 217727
rect 292671 199449 292949 199727
rect 292671 181449 292949 181727
rect 292671 163449 292949 163727
rect 292671 145449 292949 145727
rect 292671 127449 292949 127727
rect 292671 109449 292949 109727
rect 292671 91449 292949 91727
rect 292671 73449 292949 73727
rect 292671 55449 292949 55727
rect 292671 37449 292949 37727
rect 292671 19449 292949 19727
rect 292671 1449 292949 1727
rect 292671 -451 292949 -173
rect 293151 334449 293429 334727
rect 293151 316449 293429 316727
rect 293151 298449 293429 298727
rect 293151 280449 293429 280727
rect 293151 262449 293429 262727
rect 293151 244449 293429 244727
rect 293151 226449 293429 226727
rect 293151 208449 293429 208727
rect 293151 190449 293429 190727
rect 293151 172449 293429 172727
rect 293151 154449 293429 154727
rect 293151 136449 293429 136727
rect 293151 118449 293429 118727
rect 293151 100449 293429 100727
rect 293151 82449 293429 82727
rect 293151 64449 293429 64727
rect 293151 46449 293429 46727
rect 293151 28449 293429 28727
rect 293151 10449 293429 10727
rect 293151 -931 293429 -653
rect 293631 345309 293909 345587
rect 293631 327309 293909 327587
rect 293631 309309 293909 309587
rect 293631 291309 293909 291587
rect 293631 273309 293909 273587
rect 293631 255309 293909 255587
rect 293631 237309 293909 237587
rect 293631 219309 293909 219587
rect 293631 201309 293909 201587
rect 293631 183309 293909 183587
rect 293631 165309 293909 165587
rect 293631 147309 293909 147587
rect 293631 129309 293909 129587
rect 293631 111309 293909 111587
rect 293631 93309 293909 93587
rect 293631 75309 293909 75587
rect 293631 57309 293909 57587
rect 293631 39309 293909 39587
rect 293631 21309 293909 21587
rect 293631 3309 293909 3587
rect 290773 -1411 291051 -1133
rect 293631 -1411 293909 -1133
rect 294111 336309 294389 336587
rect 294111 318309 294389 318587
rect 294111 300309 294389 300587
rect 294111 282309 294389 282587
rect 294111 264309 294389 264587
rect 294111 246309 294389 246587
rect 294111 228309 294389 228587
rect 294111 210309 294389 210587
rect 294111 192309 294389 192587
rect 294111 174309 294389 174587
rect 294111 156309 294389 156587
rect 294111 138309 294389 138587
rect 294111 120309 294389 120587
rect 294111 102309 294389 102587
rect 294111 84309 294389 84587
rect 294111 66309 294389 66587
rect 294111 48309 294389 48587
rect 294111 30309 294389 30587
rect 294111 12309 294389 12587
rect 294111 -1891 294389 -1613
rect 294591 347169 294869 347447
rect 294591 329169 294869 329447
rect 294591 311169 294869 311447
rect 294591 293169 294869 293447
rect 294591 275169 294869 275447
rect 294591 257169 294869 257447
rect 294591 239169 294869 239447
rect 294591 221169 294869 221447
rect 294591 203169 294869 203447
rect 294591 185169 294869 185447
rect 294591 167169 294869 167447
rect 294591 149169 294869 149447
rect 294591 131169 294869 131447
rect 294591 113169 294869 113447
rect 294591 95169 294869 95447
rect 294591 77169 294869 77447
rect 294591 59169 294869 59447
rect 294591 41169 294869 41447
rect 294591 23169 294869 23447
rect 294591 5169 294869 5447
rect 294591 -2371 294869 -2093
rect 295071 338169 295349 338447
rect 295071 320169 295349 320447
rect 295071 302169 295349 302447
rect 295071 284169 295349 284447
rect 295071 266169 295349 266447
rect 295071 248169 295349 248447
rect 295071 230169 295349 230447
rect 295071 212169 295349 212447
rect 295071 194169 295349 194447
rect 295071 176169 295349 176447
rect 295071 158169 295349 158447
rect 295071 140169 295349 140447
rect 295071 122169 295349 122447
rect 295071 104169 295349 104447
rect 295071 86169 295349 86447
rect 295071 68169 295349 68447
rect 295071 50169 295349 50447
rect 295071 32169 295349 32447
rect 295071 14169 295349 14447
rect 295071 -2851 295349 -2573
rect 295551 349029 295829 349307
rect 295551 331029 295829 331307
rect 295551 313029 295829 313307
rect 295551 295029 295829 295307
rect 295551 277029 295829 277307
rect 295551 259029 295829 259307
rect 295551 241029 295829 241307
rect 295551 223029 295829 223307
rect 295551 205029 295829 205307
rect 295551 187029 295829 187307
rect 295551 169029 295829 169307
rect 295551 151029 295829 151307
rect 295551 133029 295829 133307
rect 295551 115029 295829 115307
rect 295551 97029 295829 97307
rect 295551 79029 295829 79307
rect 295551 61029 295829 61307
rect 295551 43029 295829 43307
rect 295551 25029 295829 25307
rect 295551 7029 295829 7307
rect 295551 -3331 295829 -3053
rect 296031 340029 296309 340307
rect 296031 322029 296309 322307
rect 296031 304029 296309 304307
rect 296031 286029 296309 286307
rect 296031 268029 296309 268307
rect 296031 250029 296309 250307
rect 296031 232029 296309 232307
rect 296031 214029 296309 214307
rect 296031 196029 296309 196307
rect 296031 178029 296309 178307
rect 296031 160029 296309 160307
rect 296031 142029 296309 142307
rect 296031 124029 296309 124307
rect 296031 106029 296309 106307
rect 296031 88029 296309 88307
rect 296031 70029 296309 70307
rect 296031 52029 296309 52307
rect 296031 34029 296309 34307
rect 296031 16029 296309 16307
rect 285493 -3811 285771 -3533
rect 296031 -3811 296309 -3533
<< metal5 >>
rect -4363 355779 296325 355795
rect -4363 355501 -4347 355779
rect -4069 355501 15493 355779
rect 15771 355501 33493 355779
rect 33771 355501 51493 355779
rect 51771 355501 69493 355779
rect 69771 355501 87493 355779
rect 87771 355501 105493 355779
rect 105771 355501 123493 355779
rect 123771 355501 141493 355779
rect 141771 355501 159493 355779
rect 159771 355501 177493 355779
rect 177771 355501 195493 355779
rect 195771 355501 213493 355779
rect 213771 355501 231493 355779
rect 231771 355501 249493 355779
rect 249771 355501 267493 355779
rect 267771 355501 285493 355779
rect 285771 355501 296031 355779
rect 296309 355501 296325 355779
rect -4363 355485 296325 355501
rect -3883 355299 295845 355315
rect -3883 355021 -3867 355299
rect -3589 355021 6493 355299
rect 6771 355021 24493 355299
rect 24771 355021 42493 355299
rect 42771 355021 60493 355299
rect 60771 355021 78493 355299
rect 78771 355021 96493 355299
rect 96771 355021 114493 355299
rect 114771 355021 132493 355299
rect 132771 355021 150493 355299
rect 150771 355021 168493 355299
rect 168771 355021 186493 355299
rect 186771 355021 204493 355299
rect 204771 355021 222493 355299
rect 222771 355021 240493 355299
rect 240771 355021 258493 355299
rect 258771 355021 276493 355299
rect 276771 355021 295551 355299
rect 295829 355021 295845 355299
rect -3883 355005 295845 355021
rect -3403 354819 295365 354835
rect -3403 354541 -3387 354819
rect -3109 354541 13633 354819
rect 13911 354541 31633 354819
rect 31911 354541 49633 354819
rect 49911 354541 67633 354819
rect 67911 354541 85633 354819
rect 85911 354541 103633 354819
rect 103911 354541 121633 354819
rect 121911 354541 139633 354819
rect 139911 354541 157633 354819
rect 157911 354541 175633 354819
rect 175911 354541 193633 354819
rect 193911 354541 211633 354819
rect 211911 354541 229633 354819
rect 229911 354541 247633 354819
rect 247911 354541 265633 354819
rect 265911 354541 283633 354819
rect 283911 354541 295071 354819
rect 295349 354541 295365 354819
rect -3403 354525 295365 354541
rect -2923 354339 294885 354355
rect -2923 354061 -2907 354339
rect -2629 354061 4633 354339
rect 4911 354061 22633 354339
rect 22911 354061 40633 354339
rect 40911 354061 58633 354339
rect 58911 354061 76633 354339
rect 76911 354061 94633 354339
rect 94911 354061 112633 354339
rect 112911 354061 130633 354339
rect 130911 354061 148633 354339
rect 148911 354061 166633 354339
rect 166911 354061 184633 354339
rect 184911 354061 202633 354339
rect 202911 354061 220633 354339
rect 220911 354061 238633 354339
rect 238911 354061 256633 354339
rect 256911 354061 274633 354339
rect 274911 354061 294591 354339
rect 294869 354061 294885 354339
rect -2923 354045 294885 354061
rect -2443 353859 294405 353875
rect -2443 353581 -2427 353859
rect -2149 353581 11773 353859
rect 12051 353581 29773 353859
rect 30051 353581 47773 353859
rect 48051 353581 65773 353859
rect 66051 353581 83773 353859
rect 84051 353581 101773 353859
rect 102051 353581 119773 353859
rect 120051 353581 137773 353859
rect 138051 353581 155773 353859
rect 156051 353581 173773 353859
rect 174051 353581 191773 353859
rect 192051 353581 209773 353859
rect 210051 353581 227773 353859
rect 228051 353581 245773 353859
rect 246051 353581 263773 353859
rect 264051 353581 281773 353859
rect 282051 353581 294111 353859
rect 294389 353581 294405 353859
rect -2443 353565 294405 353581
rect -1963 353379 293925 353395
rect -1963 353101 -1947 353379
rect -1669 353101 2773 353379
rect 3051 353101 20773 353379
rect 21051 353101 38773 353379
rect 39051 353101 56773 353379
rect 57051 353101 74773 353379
rect 75051 353101 92773 353379
rect 93051 353101 110773 353379
rect 111051 353101 128773 353379
rect 129051 353101 146773 353379
rect 147051 353101 164773 353379
rect 165051 353101 182773 353379
rect 183051 353101 200773 353379
rect 201051 353101 218773 353379
rect 219051 353101 236773 353379
rect 237051 353101 254773 353379
rect 255051 353101 272773 353379
rect 273051 353101 290773 353379
rect 291051 353101 293631 353379
rect 293909 353101 293925 353379
rect -1963 353085 293925 353101
rect -1483 352899 293445 352915
rect -1483 352621 -1467 352899
rect -1189 352621 9913 352899
rect 10191 352621 27913 352899
rect 28191 352621 45913 352899
rect 46191 352621 63913 352899
rect 64191 352621 81913 352899
rect 82191 352621 99913 352899
rect 100191 352621 117913 352899
rect 118191 352621 135913 352899
rect 136191 352621 153913 352899
rect 154191 352621 171913 352899
rect 172191 352621 189913 352899
rect 190191 352621 207913 352899
rect 208191 352621 225913 352899
rect 226191 352621 243913 352899
rect 244191 352621 261913 352899
rect 262191 352621 279913 352899
rect 280191 352621 293151 352899
rect 293429 352621 293445 352899
rect -1483 352605 293445 352621
rect -1003 352419 292965 352435
rect -1003 352141 -987 352419
rect -709 352141 913 352419
rect 1191 352141 18913 352419
rect 19191 352141 36913 352419
rect 37191 352141 54913 352419
rect 55191 352141 72913 352419
rect 73191 352141 90913 352419
rect 91191 352141 108913 352419
rect 109191 352141 126913 352419
rect 127191 352141 144913 352419
rect 145191 352141 162913 352419
rect 163191 352141 180913 352419
rect 181191 352141 198913 352419
rect 199191 352141 216913 352419
rect 217191 352141 234913 352419
rect 235191 352141 252913 352419
rect 253191 352141 270913 352419
rect 271191 352141 288913 352419
rect 289191 352141 292671 352419
rect 292949 352141 292965 352419
rect -1003 352125 292965 352141
rect -4363 349307 296325 349323
rect -4363 349029 -3867 349307
rect -3589 349029 6493 349307
rect 6771 349029 24493 349307
rect 24771 349029 42493 349307
rect 42771 349029 60493 349307
rect 60771 349029 78493 349307
rect 78771 349029 96493 349307
rect 96771 349029 114493 349307
rect 114771 349029 132493 349307
rect 132771 349029 150493 349307
rect 150771 349029 168493 349307
rect 168771 349029 186493 349307
rect 186771 349029 204493 349307
rect 204771 349029 222493 349307
rect 222771 349029 240493 349307
rect 240771 349029 258493 349307
rect 258771 349029 276493 349307
rect 276771 349029 295551 349307
rect 295829 349029 296325 349307
rect -4363 349013 296325 349029
rect -3403 347447 295365 347463
rect -3403 347169 -2907 347447
rect -2629 347169 4633 347447
rect 4911 347169 22633 347447
rect 22911 347169 40633 347447
rect 40911 347169 58633 347447
rect 58911 347169 76633 347447
rect 76911 347169 94633 347447
rect 94911 347169 112633 347447
rect 112911 347169 130633 347447
rect 130911 347169 148633 347447
rect 148911 347169 166633 347447
rect 166911 347169 184633 347447
rect 184911 347169 202633 347447
rect 202911 347169 220633 347447
rect 220911 347169 238633 347447
rect 238911 347169 256633 347447
rect 256911 347169 274633 347447
rect 274911 347169 294591 347447
rect 294869 347169 295365 347447
rect -3403 347153 295365 347169
rect -2443 345587 294405 345603
rect -2443 345309 -1947 345587
rect -1669 345309 2773 345587
rect 3051 345309 20773 345587
rect 21051 345309 38773 345587
rect 39051 345309 56773 345587
rect 57051 345309 74773 345587
rect 75051 345309 92773 345587
rect 93051 345309 110773 345587
rect 111051 345309 128773 345587
rect 129051 345309 146773 345587
rect 147051 345309 164773 345587
rect 165051 345309 182773 345587
rect 183051 345309 200773 345587
rect 201051 345309 218773 345587
rect 219051 345309 236773 345587
rect 237051 345309 254773 345587
rect 255051 345309 272773 345587
rect 273051 345309 290773 345587
rect 291051 345309 293631 345587
rect 293909 345309 294405 345587
rect -2443 345293 294405 345309
rect -1483 343727 293445 343743
rect -1483 343449 -987 343727
rect -709 343449 913 343727
rect 1191 343449 18913 343727
rect 19191 343449 36913 343727
rect 37191 343449 54913 343727
rect 55191 343449 72913 343727
rect 73191 343449 90913 343727
rect 91191 343449 108913 343727
rect 109191 343449 126913 343727
rect 127191 343449 144913 343727
rect 145191 343449 162913 343727
rect 163191 343449 180913 343727
rect 181191 343449 198913 343727
rect 199191 343449 216913 343727
rect 217191 343449 234913 343727
rect 235191 343449 252913 343727
rect 253191 343449 270913 343727
rect 271191 343449 288913 343727
rect 289191 343449 292671 343727
rect 292949 343449 293445 343727
rect -1483 343433 293445 343449
rect -4363 340307 296325 340323
rect -4363 340029 -4347 340307
rect -4069 340029 15493 340307
rect 15771 340029 33493 340307
rect 33771 340029 51493 340307
rect 51771 340029 69493 340307
rect 69771 340029 87493 340307
rect 87771 340029 105493 340307
rect 105771 340029 123493 340307
rect 123771 340029 141493 340307
rect 141771 340029 159493 340307
rect 159771 340029 177493 340307
rect 177771 340029 195493 340307
rect 195771 340029 213493 340307
rect 213771 340029 231493 340307
rect 231771 340029 249493 340307
rect 249771 340029 267493 340307
rect 267771 340029 285493 340307
rect 285771 340029 296031 340307
rect 296309 340029 296325 340307
rect -4363 340013 296325 340029
rect -3403 338447 295365 338463
rect -3403 338169 -3387 338447
rect -3109 338169 13633 338447
rect 13911 338169 31633 338447
rect 31911 338169 49633 338447
rect 49911 338169 67633 338447
rect 67911 338169 85633 338447
rect 85911 338169 103633 338447
rect 103911 338169 121633 338447
rect 121911 338169 139633 338447
rect 139911 338169 157633 338447
rect 157911 338169 175633 338447
rect 175911 338169 193633 338447
rect 193911 338169 211633 338447
rect 211911 338169 229633 338447
rect 229911 338169 247633 338447
rect 247911 338169 265633 338447
rect 265911 338169 283633 338447
rect 283911 338169 295071 338447
rect 295349 338169 295365 338447
rect -3403 338153 295365 338169
rect -2443 336587 294405 336603
rect -2443 336309 -2427 336587
rect -2149 336309 11773 336587
rect 12051 336309 29773 336587
rect 30051 336309 47773 336587
rect 48051 336309 65773 336587
rect 66051 336309 83773 336587
rect 84051 336309 101773 336587
rect 102051 336309 119773 336587
rect 120051 336309 137773 336587
rect 138051 336309 155773 336587
rect 156051 336309 173773 336587
rect 174051 336309 191773 336587
rect 192051 336309 209773 336587
rect 210051 336309 227773 336587
rect 228051 336309 245773 336587
rect 246051 336309 263773 336587
rect 264051 336309 281773 336587
rect 282051 336309 294111 336587
rect 294389 336309 294405 336587
rect -2443 336293 294405 336309
rect -1483 334727 293445 334743
rect -1483 334449 -1467 334727
rect -1189 334449 9913 334727
rect 10191 334449 27913 334727
rect 28191 334449 45913 334727
rect 46191 334449 63913 334727
rect 64191 334449 81913 334727
rect 82191 334449 99913 334727
rect 100191 334449 117913 334727
rect 118191 334449 135913 334727
rect 136191 334449 153913 334727
rect 154191 334449 171913 334727
rect 172191 334449 189913 334727
rect 190191 334449 207913 334727
rect 208191 334449 225913 334727
rect 226191 334449 243913 334727
rect 244191 334449 261913 334727
rect 262191 334449 279913 334727
rect 280191 334449 293151 334727
rect 293429 334449 293445 334727
rect -1483 334433 293445 334449
rect -4363 331307 296325 331323
rect -4363 331029 -3867 331307
rect -3589 331029 6493 331307
rect 6771 331029 24493 331307
rect 24771 331029 42493 331307
rect 42771 331029 60493 331307
rect 60771 331029 78493 331307
rect 78771 331029 96493 331307
rect 96771 331029 114493 331307
rect 114771 331029 132493 331307
rect 132771 331029 150493 331307
rect 150771 331029 168493 331307
rect 168771 331029 186493 331307
rect 186771 331029 204493 331307
rect 204771 331029 222493 331307
rect 222771 331029 240493 331307
rect 240771 331029 258493 331307
rect 258771 331029 276493 331307
rect 276771 331029 295551 331307
rect 295829 331029 296325 331307
rect -4363 331013 296325 331029
rect -3403 329447 295365 329463
rect -3403 329169 -2907 329447
rect -2629 329169 4633 329447
rect 4911 329169 22633 329447
rect 22911 329169 40633 329447
rect 40911 329169 58633 329447
rect 58911 329169 76633 329447
rect 76911 329169 94633 329447
rect 94911 329169 112633 329447
rect 112911 329169 130633 329447
rect 130911 329169 148633 329447
rect 148911 329169 166633 329447
rect 166911 329169 184633 329447
rect 184911 329169 202633 329447
rect 202911 329169 220633 329447
rect 220911 329169 238633 329447
rect 238911 329169 256633 329447
rect 256911 329169 274633 329447
rect 274911 329169 294591 329447
rect 294869 329169 295365 329447
rect -3403 329153 295365 329169
rect -2443 327587 294405 327603
rect -2443 327309 -1947 327587
rect -1669 327309 2773 327587
rect 3051 327309 20773 327587
rect 21051 327309 38773 327587
rect 39051 327309 56773 327587
rect 57051 327309 74773 327587
rect 75051 327309 92773 327587
rect 93051 327309 110773 327587
rect 111051 327309 128773 327587
rect 129051 327309 146773 327587
rect 147051 327309 164773 327587
rect 165051 327309 182773 327587
rect 183051 327309 200773 327587
rect 201051 327309 218773 327587
rect 219051 327309 236773 327587
rect 237051 327309 254773 327587
rect 255051 327309 272773 327587
rect 273051 327309 290773 327587
rect 291051 327309 293631 327587
rect 293909 327309 294405 327587
rect -2443 327293 294405 327309
rect -1483 325727 293445 325743
rect -1483 325449 -987 325727
rect -709 325449 913 325727
rect 1191 325449 18913 325727
rect 19191 325449 36913 325727
rect 37191 325449 54913 325727
rect 55191 325449 72913 325727
rect 73191 325449 90913 325727
rect 91191 325449 108913 325727
rect 109191 325449 126913 325727
rect 127191 325449 144913 325727
rect 145191 325449 162913 325727
rect 163191 325449 180913 325727
rect 181191 325449 198913 325727
rect 199191 325449 216913 325727
rect 217191 325449 234913 325727
rect 235191 325449 252913 325727
rect 253191 325449 270913 325727
rect 271191 325449 288913 325727
rect 289191 325449 292671 325727
rect 292949 325449 293445 325727
rect -1483 325433 293445 325449
rect -4363 322307 296325 322323
rect -4363 322029 -4347 322307
rect -4069 322029 15493 322307
rect 15771 322029 33493 322307
rect 33771 322029 51493 322307
rect 51771 322029 69493 322307
rect 69771 322029 87493 322307
rect 87771 322029 105493 322307
rect 105771 322029 123493 322307
rect 123771 322029 141493 322307
rect 141771 322029 159493 322307
rect 159771 322029 177493 322307
rect 177771 322029 195493 322307
rect 195771 322029 213493 322307
rect 213771 322029 231493 322307
rect 231771 322029 249493 322307
rect 249771 322029 267493 322307
rect 267771 322029 285493 322307
rect 285771 322029 296031 322307
rect 296309 322029 296325 322307
rect -4363 322013 296325 322029
rect -3403 320447 295365 320463
rect -3403 320169 -3387 320447
rect -3109 320169 13633 320447
rect 13911 320169 31633 320447
rect 31911 320169 49633 320447
rect 49911 320169 67633 320447
rect 67911 320169 85633 320447
rect 85911 320169 103633 320447
rect 103911 320169 121633 320447
rect 121911 320169 139633 320447
rect 139911 320169 157633 320447
rect 157911 320169 175633 320447
rect 175911 320169 193633 320447
rect 193911 320169 211633 320447
rect 211911 320169 229633 320447
rect 229911 320169 247633 320447
rect 247911 320169 265633 320447
rect 265911 320169 283633 320447
rect 283911 320169 295071 320447
rect 295349 320169 295365 320447
rect -3403 320153 295365 320169
rect -2443 318587 294405 318603
rect -2443 318309 -2427 318587
rect -2149 318309 11773 318587
rect 12051 318309 29773 318587
rect 30051 318309 47773 318587
rect 48051 318309 65773 318587
rect 66051 318309 83773 318587
rect 84051 318309 101773 318587
rect 102051 318309 119773 318587
rect 120051 318309 137773 318587
rect 138051 318309 155773 318587
rect 156051 318309 173773 318587
rect 174051 318309 191773 318587
rect 192051 318309 209773 318587
rect 210051 318309 227773 318587
rect 228051 318309 245773 318587
rect 246051 318309 263773 318587
rect 264051 318309 281773 318587
rect 282051 318309 294111 318587
rect 294389 318309 294405 318587
rect -2443 318293 294405 318309
rect -1483 316727 293445 316743
rect -1483 316449 -1467 316727
rect -1189 316449 9913 316727
rect 10191 316449 27913 316727
rect 28191 316449 45913 316727
rect 46191 316449 63913 316727
rect 64191 316449 81913 316727
rect 82191 316449 99913 316727
rect 100191 316449 117913 316727
rect 118191 316449 135913 316727
rect 136191 316449 153913 316727
rect 154191 316449 171913 316727
rect 172191 316449 189913 316727
rect 190191 316449 207913 316727
rect 208191 316449 225913 316727
rect 226191 316449 243913 316727
rect 244191 316449 261913 316727
rect 262191 316449 279913 316727
rect 280191 316449 293151 316727
rect 293429 316449 293445 316727
rect -1483 316433 293445 316449
rect -4363 313307 296325 313323
rect -4363 313029 -3867 313307
rect -3589 313029 6493 313307
rect 6771 313029 24493 313307
rect 24771 313029 42493 313307
rect 42771 313029 60493 313307
rect 60771 313029 78493 313307
rect 78771 313029 96493 313307
rect 96771 313029 114493 313307
rect 114771 313029 132493 313307
rect 132771 313029 150493 313307
rect 150771 313029 168493 313307
rect 168771 313029 186493 313307
rect 186771 313029 204493 313307
rect 204771 313029 222493 313307
rect 222771 313029 240493 313307
rect 240771 313029 258493 313307
rect 258771 313029 276493 313307
rect 276771 313029 295551 313307
rect 295829 313029 296325 313307
rect -4363 313013 296325 313029
rect -3403 311447 295365 311463
rect -3403 311169 -2907 311447
rect -2629 311169 4633 311447
rect 4911 311169 22633 311447
rect 22911 311169 40633 311447
rect 40911 311169 58633 311447
rect 58911 311169 76633 311447
rect 76911 311169 94633 311447
rect 94911 311169 112633 311447
rect 112911 311169 130633 311447
rect 130911 311169 148633 311447
rect 148911 311169 166633 311447
rect 166911 311169 184633 311447
rect 184911 311169 202633 311447
rect 202911 311169 220633 311447
rect 220911 311169 238633 311447
rect 238911 311169 256633 311447
rect 256911 311169 274633 311447
rect 274911 311169 294591 311447
rect 294869 311169 295365 311447
rect -3403 311153 295365 311169
rect -2443 309587 294405 309603
rect -2443 309309 -1947 309587
rect -1669 309309 2773 309587
rect 3051 309309 20773 309587
rect 21051 309309 38773 309587
rect 39051 309309 56773 309587
rect 57051 309309 74773 309587
rect 75051 309309 92773 309587
rect 93051 309309 110773 309587
rect 111051 309309 128773 309587
rect 129051 309309 146773 309587
rect 147051 309309 164773 309587
rect 165051 309309 182773 309587
rect 183051 309309 200773 309587
rect 201051 309309 218773 309587
rect 219051 309309 236773 309587
rect 237051 309309 254773 309587
rect 255051 309309 272773 309587
rect 273051 309309 290773 309587
rect 291051 309309 293631 309587
rect 293909 309309 294405 309587
rect -2443 309293 294405 309309
rect -1483 307727 293445 307743
rect -1483 307449 -987 307727
rect -709 307449 913 307727
rect 1191 307449 18913 307727
rect 19191 307449 36913 307727
rect 37191 307449 54913 307727
rect 55191 307449 72913 307727
rect 73191 307449 90913 307727
rect 91191 307449 108913 307727
rect 109191 307449 126913 307727
rect 127191 307449 144913 307727
rect 145191 307449 162913 307727
rect 163191 307449 180913 307727
rect 181191 307449 198913 307727
rect 199191 307449 216913 307727
rect 217191 307449 234913 307727
rect 235191 307449 252913 307727
rect 253191 307449 270913 307727
rect 271191 307449 288913 307727
rect 289191 307449 292671 307727
rect 292949 307449 293445 307727
rect -1483 307433 293445 307449
rect -4363 304307 296325 304323
rect -4363 304029 -4347 304307
rect -4069 304029 15493 304307
rect 15771 304029 33493 304307
rect 33771 304029 51493 304307
rect 51771 304029 69493 304307
rect 69771 304029 87493 304307
rect 87771 304029 105493 304307
rect 105771 304029 123493 304307
rect 123771 304029 141493 304307
rect 141771 304029 159493 304307
rect 159771 304029 177493 304307
rect 177771 304029 195493 304307
rect 195771 304029 213493 304307
rect 213771 304029 231493 304307
rect 231771 304029 249493 304307
rect 249771 304029 267493 304307
rect 267771 304029 285493 304307
rect 285771 304029 296031 304307
rect 296309 304029 296325 304307
rect -4363 304013 296325 304029
rect -3403 302447 295365 302463
rect -3403 302169 -3387 302447
rect -3109 302169 13633 302447
rect 13911 302169 31633 302447
rect 31911 302169 49633 302447
rect 49911 302169 67633 302447
rect 67911 302169 85633 302447
rect 85911 302169 103633 302447
rect 103911 302169 121633 302447
rect 121911 302169 139633 302447
rect 139911 302169 157633 302447
rect 157911 302169 175633 302447
rect 175911 302169 193633 302447
rect 193911 302169 211633 302447
rect 211911 302169 229633 302447
rect 229911 302169 247633 302447
rect 247911 302169 265633 302447
rect 265911 302169 283633 302447
rect 283911 302169 295071 302447
rect 295349 302169 295365 302447
rect -3403 302153 295365 302169
rect -2443 300587 294405 300603
rect -2443 300309 -2427 300587
rect -2149 300309 11773 300587
rect 12051 300309 29773 300587
rect 30051 300309 47773 300587
rect 48051 300309 65773 300587
rect 66051 300309 83773 300587
rect 84051 300309 101773 300587
rect 102051 300309 119773 300587
rect 120051 300309 137773 300587
rect 138051 300309 155773 300587
rect 156051 300309 173773 300587
rect 174051 300309 191773 300587
rect 192051 300309 209773 300587
rect 210051 300309 227773 300587
rect 228051 300309 245773 300587
rect 246051 300309 263773 300587
rect 264051 300309 281773 300587
rect 282051 300309 294111 300587
rect 294389 300309 294405 300587
rect -2443 300293 294405 300309
rect -1483 298727 293445 298743
rect -1483 298449 -1467 298727
rect -1189 298449 9913 298727
rect 10191 298449 27913 298727
rect 28191 298449 45913 298727
rect 46191 298449 63913 298727
rect 64191 298449 81913 298727
rect 82191 298449 99913 298727
rect 100191 298449 117913 298727
rect 118191 298449 135913 298727
rect 136191 298449 153913 298727
rect 154191 298449 171913 298727
rect 172191 298449 189913 298727
rect 190191 298449 207913 298727
rect 208191 298449 225913 298727
rect 226191 298449 243913 298727
rect 244191 298449 261913 298727
rect 262191 298449 279913 298727
rect 280191 298449 293151 298727
rect 293429 298449 293445 298727
rect -1483 298433 293445 298449
rect -4363 295307 296325 295323
rect -4363 295029 -3867 295307
rect -3589 295029 6493 295307
rect 6771 295029 24493 295307
rect 24771 295029 42493 295307
rect 42771 295029 60493 295307
rect 60771 295029 78493 295307
rect 78771 295029 96493 295307
rect 96771 295029 114493 295307
rect 114771 295029 132493 295307
rect 132771 295029 150493 295307
rect 150771 295029 168493 295307
rect 168771 295029 186493 295307
rect 186771 295029 204493 295307
rect 204771 295029 222493 295307
rect 222771 295029 240493 295307
rect 240771 295029 258493 295307
rect 258771 295029 276493 295307
rect 276771 295029 295551 295307
rect 295829 295029 296325 295307
rect -4363 295013 296325 295029
rect -3403 293447 295365 293463
rect -3403 293169 -2907 293447
rect -2629 293169 4633 293447
rect 4911 293169 22633 293447
rect 22911 293169 40633 293447
rect 40911 293169 58633 293447
rect 58911 293169 76633 293447
rect 76911 293169 94633 293447
rect 94911 293169 112633 293447
rect 112911 293169 130633 293447
rect 130911 293169 148633 293447
rect 148911 293169 166633 293447
rect 166911 293169 184633 293447
rect 184911 293169 202633 293447
rect 202911 293169 220633 293447
rect 220911 293169 238633 293447
rect 238911 293169 256633 293447
rect 256911 293169 274633 293447
rect 274911 293169 294591 293447
rect 294869 293169 295365 293447
rect -3403 293153 295365 293169
rect -2443 291587 294405 291603
rect -2443 291309 -1947 291587
rect -1669 291309 2773 291587
rect 3051 291309 20773 291587
rect 21051 291309 38773 291587
rect 39051 291309 56773 291587
rect 57051 291309 74773 291587
rect 75051 291309 92773 291587
rect 93051 291309 110773 291587
rect 111051 291309 128773 291587
rect 129051 291309 146773 291587
rect 147051 291309 164773 291587
rect 165051 291309 182773 291587
rect 183051 291309 200773 291587
rect 201051 291309 218773 291587
rect 219051 291309 236773 291587
rect 237051 291309 254773 291587
rect 255051 291309 272773 291587
rect 273051 291309 290773 291587
rect 291051 291309 293631 291587
rect 293909 291309 294405 291587
rect -2443 291293 294405 291309
rect -1483 289727 293445 289743
rect -1483 289449 -987 289727
rect -709 289449 913 289727
rect 1191 289449 18913 289727
rect 19191 289449 36913 289727
rect 37191 289449 54913 289727
rect 55191 289449 72913 289727
rect 73191 289449 90913 289727
rect 91191 289449 108913 289727
rect 109191 289449 126913 289727
rect 127191 289449 144913 289727
rect 145191 289449 162913 289727
rect 163191 289449 180913 289727
rect 181191 289449 198913 289727
rect 199191 289449 216913 289727
rect 217191 289449 234913 289727
rect 235191 289449 252913 289727
rect 253191 289449 270913 289727
rect 271191 289449 288913 289727
rect 289191 289449 292671 289727
rect 292949 289449 293445 289727
rect -1483 289433 293445 289449
rect -4363 286307 296325 286323
rect -4363 286029 -4347 286307
rect -4069 286029 15493 286307
rect 15771 286029 33493 286307
rect 33771 286029 51493 286307
rect 51771 286029 69493 286307
rect 69771 286029 87493 286307
rect 87771 286029 105493 286307
rect 105771 286029 123493 286307
rect 123771 286029 141493 286307
rect 141771 286029 159493 286307
rect 159771 286029 177493 286307
rect 177771 286029 195493 286307
rect 195771 286029 213493 286307
rect 213771 286029 231493 286307
rect 231771 286029 249493 286307
rect 249771 286029 267493 286307
rect 267771 286029 285493 286307
rect 285771 286029 296031 286307
rect 296309 286029 296325 286307
rect -4363 286013 296325 286029
rect -3403 284447 295365 284463
rect -3403 284169 -3387 284447
rect -3109 284169 13633 284447
rect 13911 284169 31633 284447
rect 31911 284169 49633 284447
rect 49911 284169 67633 284447
rect 67911 284169 85633 284447
rect 85911 284169 103633 284447
rect 103911 284169 121633 284447
rect 121911 284169 139633 284447
rect 139911 284169 157633 284447
rect 157911 284169 175633 284447
rect 175911 284169 193633 284447
rect 193911 284169 211633 284447
rect 211911 284169 229633 284447
rect 229911 284169 247633 284447
rect 247911 284169 265633 284447
rect 265911 284169 283633 284447
rect 283911 284169 295071 284447
rect 295349 284169 295365 284447
rect -3403 284153 295365 284169
rect -2443 282587 294405 282603
rect -2443 282309 -2427 282587
rect -2149 282309 11773 282587
rect 12051 282309 29773 282587
rect 30051 282309 47773 282587
rect 48051 282309 65773 282587
rect 66051 282309 83773 282587
rect 84051 282309 101773 282587
rect 102051 282309 119773 282587
rect 120051 282309 137773 282587
rect 138051 282309 155773 282587
rect 156051 282309 173773 282587
rect 174051 282309 191773 282587
rect 192051 282309 209773 282587
rect 210051 282309 227773 282587
rect 228051 282309 245773 282587
rect 246051 282309 263773 282587
rect 264051 282309 281773 282587
rect 282051 282309 294111 282587
rect 294389 282309 294405 282587
rect -2443 282293 294405 282309
rect -1483 280727 293445 280743
rect -1483 280449 -1467 280727
rect -1189 280449 9913 280727
rect 10191 280449 27913 280727
rect 28191 280449 45913 280727
rect 46191 280449 63913 280727
rect 64191 280449 81913 280727
rect 82191 280449 99913 280727
rect 100191 280449 117913 280727
rect 118191 280449 135913 280727
rect 136191 280449 153913 280727
rect 154191 280449 171913 280727
rect 172191 280449 189913 280727
rect 190191 280449 207913 280727
rect 208191 280449 225913 280727
rect 226191 280449 243913 280727
rect 244191 280449 261913 280727
rect 262191 280449 279913 280727
rect 280191 280449 293151 280727
rect 293429 280449 293445 280727
rect -1483 280433 293445 280449
rect -4363 277307 296325 277323
rect -4363 277029 -3867 277307
rect -3589 277029 6493 277307
rect 6771 277029 24493 277307
rect 24771 277029 42493 277307
rect 42771 277029 60493 277307
rect 60771 277029 78493 277307
rect 78771 277029 96493 277307
rect 96771 277029 114493 277307
rect 114771 277029 132493 277307
rect 132771 277029 150493 277307
rect 150771 277029 168493 277307
rect 168771 277029 186493 277307
rect 186771 277029 204493 277307
rect 204771 277029 222493 277307
rect 222771 277029 240493 277307
rect 240771 277029 258493 277307
rect 258771 277029 276493 277307
rect 276771 277029 295551 277307
rect 295829 277029 296325 277307
rect -4363 277013 296325 277029
rect -3403 275447 295365 275463
rect -3403 275169 -2907 275447
rect -2629 275169 4633 275447
rect 4911 275169 22633 275447
rect 22911 275169 40633 275447
rect 40911 275169 58633 275447
rect 58911 275169 76633 275447
rect 76911 275169 94633 275447
rect 94911 275169 112633 275447
rect 112911 275169 130633 275447
rect 130911 275169 148633 275447
rect 148911 275169 166633 275447
rect 166911 275169 184633 275447
rect 184911 275169 202633 275447
rect 202911 275169 220633 275447
rect 220911 275169 238633 275447
rect 238911 275169 256633 275447
rect 256911 275169 274633 275447
rect 274911 275169 294591 275447
rect 294869 275169 295365 275447
rect -3403 275153 295365 275169
rect -2443 273587 294405 273603
rect -2443 273309 -1947 273587
rect -1669 273309 2773 273587
rect 3051 273309 20773 273587
rect 21051 273309 38773 273587
rect 39051 273309 56773 273587
rect 57051 273309 74773 273587
rect 75051 273309 92773 273587
rect 93051 273309 110773 273587
rect 111051 273309 128773 273587
rect 129051 273309 146773 273587
rect 147051 273309 164773 273587
rect 165051 273309 182773 273587
rect 183051 273309 200773 273587
rect 201051 273309 218773 273587
rect 219051 273309 236773 273587
rect 237051 273309 254773 273587
rect 255051 273309 272773 273587
rect 273051 273309 290773 273587
rect 291051 273309 293631 273587
rect 293909 273309 294405 273587
rect -2443 273293 294405 273309
rect -1483 271727 293445 271743
rect -1483 271449 -987 271727
rect -709 271449 913 271727
rect 1191 271449 18913 271727
rect 19191 271449 36913 271727
rect 37191 271449 54913 271727
rect 55191 271449 72913 271727
rect 73191 271449 90913 271727
rect 91191 271449 108913 271727
rect 109191 271449 126913 271727
rect 127191 271449 144913 271727
rect 145191 271449 162913 271727
rect 163191 271449 180913 271727
rect 181191 271449 198913 271727
rect 199191 271449 216913 271727
rect 217191 271449 234913 271727
rect 235191 271449 252913 271727
rect 253191 271449 270913 271727
rect 271191 271449 288913 271727
rect 289191 271449 292671 271727
rect 292949 271449 293445 271727
rect -1483 271433 293445 271449
rect -4363 268307 296325 268323
rect -4363 268029 -4347 268307
rect -4069 268029 15493 268307
rect 15771 268029 33493 268307
rect 33771 268029 51493 268307
rect 51771 268029 69493 268307
rect 69771 268029 87493 268307
rect 87771 268029 105493 268307
rect 105771 268029 123493 268307
rect 123771 268029 141493 268307
rect 141771 268029 159493 268307
rect 159771 268029 177493 268307
rect 177771 268029 195493 268307
rect 195771 268029 213493 268307
rect 213771 268029 231493 268307
rect 231771 268029 249493 268307
rect 249771 268029 267493 268307
rect 267771 268029 285493 268307
rect 285771 268029 296031 268307
rect 296309 268029 296325 268307
rect -4363 268013 296325 268029
rect -3403 266447 295365 266463
rect -3403 266169 -3387 266447
rect -3109 266169 13633 266447
rect 13911 266169 31633 266447
rect 31911 266169 49633 266447
rect 49911 266169 67633 266447
rect 67911 266169 85633 266447
rect 85911 266169 103633 266447
rect 103911 266169 121633 266447
rect 121911 266169 139633 266447
rect 139911 266169 157633 266447
rect 157911 266169 175633 266447
rect 175911 266169 193633 266447
rect 193911 266169 211633 266447
rect 211911 266169 229633 266447
rect 229911 266169 247633 266447
rect 247911 266169 265633 266447
rect 265911 266169 283633 266447
rect 283911 266169 295071 266447
rect 295349 266169 295365 266447
rect -3403 266153 295365 266169
rect -2443 264587 294405 264603
rect -2443 264309 -2427 264587
rect -2149 264309 11773 264587
rect 12051 264309 29773 264587
rect 30051 264309 47773 264587
rect 48051 264309 65773 264587
rect 66051 264309 83773 264587
rect 84051 264309 101773 264587
rect 102051 264309 119773 264587
rect 120051 264309 137773 264587
rect 138051 264309 155773 264587
rect 156051 264309 173773 264587
rect 174051 264309 191773 264587
rect 192051 264309 209773 264587
rect 210051 264309 227773 264587
rect 228051 264309 245773 264587
rect 246051 264309 263773 264587
rect 264051 264309 281773 264587
rect 282051 264309 294111 264587
rect 294389 264309 294405 264587
rect -2443 264293 294405 264309
rect -1483 262727 293445 262743
rect -1483 262449 -1467 262727
rect -1189 262449 9913 262727
rect 10191 262449 27913 262727
rect 28191 262449 45913 262727
rect 46191 262449 63913 262727
rect 64191 262449 81913 262727
rect 82191 262449 99913 262727
rect 100191 262449 117913 262727
rect 118191 262449 135913 262727
rect 136191 262449 153913 262727
rect 154191 262449 171913 262727
rect 172191 262449 189913 262727
rect 190191 262449 207913 262727
rect 208191 262449 225913 262727
rect 226191 262449 243913 262727
rect 244191 262449 261913 262727
rect 262191 262449 279913 262727
rect 280191 262449 293151 262727
rect 293429 262449 293445 262727
rect -1483 262433 293445 262449
rect -4363 259307 296325 259323
rect -4363 259029 -3867 259307
rect -3589 259029 6493 259307
rect 6771 259029 24493 259307
rect 24771 259029 42493 259307
rect 42771 259029 60493 259307
rect 60771 259029 78493 259307
rect 78771 259029 96493 259307
rect 96771 259029 114493 259307
rect 114771 259029 132493 259307
rect 132771 259029 150493 259307
rect 150771 259029 168493 259307
rect 168771 259029 186493 259307
rect 186771 259029 204493 259307
rect 204771 259029 222493 259307
rect 222771 259029 240493 259307
rect 240771 259029 258493 259307
rect 258771 259029 276493 259307
rect 276771 259029 295551 259307
rect 295829 259029 296325 259307
rect -4363 259013 296325 259029
rect -3403 257447 295365 257463
rect -3403 257169 -2907 257447
rect -2629 257169 4633 257447
rect 4911 257169 22633 257447
rect 22911 257169 40633 257447
rect 40911 257169 58633 257447
rect 58911 257169 76633 257447
rect 76911 257169 94633 257447
rect 94911 257169 112633 257447
rect 112911 257169 130633 257447
rect 130911 257169 148633 257447
rect 148911 257169 166633 257447
rect 166911 257169 184633 257447
rect 184911 257169 202633 257447
rect 202911 257169 220633 257447
rect 220911 257169 238633 257447
rect 238911 257169 256633 257447
rect 256911 257169 274633 257447
rect 274911 257169 294591 257447
rect 294869 257169 295365 257447
rect -3403 257153 295365 257169
rect -2443 255587 294405 255603
rect -2443 255309 -1947 255587
rect -1669 255309 2773 255587
rect 3051 255309 20773 255587
rect 21051 255309 38773 255587
rect 39051 255309 56773 255587
rect 57051 255309 74773 255587
rect 75051 255309 92773 255587
rect 93051 255309 110773 255587
rect 111051 255309 128773 255587
rect 129051 255309 146773 255587
rect 147051 255309 164773 255587
rect 165051 255309 182773 255587
rect 183051 255309 200773 255587
rect 201051 255309 218773 255587
rect 219051 255309 236773 255587
rect 237051 255309 254773 255587
rect 255051 255309 272773 255587
rect 273051 255309 290773 255587
rect 291051 255309 293631 255587
rect 293909 255309 294405 255587
rect -2443 255293 294405 255309
rect -1483 253727 293445 253743
rect -1483 253449 -987 253727
rect -709 253449 913 253727
rect 1191 253449 18913 253727
rect 19191 253449 36913 253727
rect 37191 253449 54913 253727
rect 55191 253449 72913 253727
rect 73191 253449 90913 253727
rect 91191 253449 108913 253727
rect 109191 253449 126913 253727
rect 127191 253449 144913 253727
rect 145191 253449 162913 253727
rect 163191 253449 180913 253727
rect 181191 253449 198913 253727
rect 199191 253449 216913 253727
rect 217191 253449 234913 253727
rect 235191 253449 252913 253727
rect 253191 253449 270913 253727
rect 271191 253449 288913 253727
rect 289191 253449 292671 253727
rect 292949 253449 293445 253727
rect -1483 253433 293445 253449
rect -4363 250307 296325 250323
rect -4363 250029 -4347 250307
rect -4069 250029 15493 250307
rect 15771 250029 33493 250307
rect 33771 250029 51493 250307
rect 51771 250029 69493 250307
rect 69771 250029 87493 250307
rect 87771 250029 105493 250307
rect 105771 250029 123493 250307
rect 123771 250029 141493 250307
rect 141771 250029 159493 250307
rect 159771 250029 177493 250307
rect 177771 250029 195493 250307
rect 195771 250029 213493 250307
rect 213771 250029 231493 250307
rect 231771 250029 249493 250307
rect 249771 250029 267493 250307
rect 267771 250029 285493 250307
rect 285771 250029 296031 250307
rect 296309 250029 296325 250307
rect -4363 250013 296325 250029
rect -3403 248447 295365 248463
rect -3403 248169 -3387 248447
rect -3109 248169 13633 248447
rect 13911 248169 31633 248447
rect 31911 248169 49633 248447
rect 49911 248169 67633 248447
rect 67911 248169 85633 248447
rect 85911 248169 103633 248447
rect 103911 248169 121633 248447
rect 121911 248169 139633 248447
rect 139911 248169 157633 248447
rect 157911 248169 175633 248447
rect 175911 248169 193633 248447
rect 193911 248169 211633 248447
rect 211911 248169 229633 248447
rect 229911 248169 247633 248447
rect 247911 248169 265633 248447
rect 265911 248169 283633 248447
rect 283911 248169 295071 248447
rect 295349 248169 295365 248447
rect -3403 248153 295365 248169
rect -2443 246587 294405 246603
rect -2443 246309 -2427 246587
rect -2149 246309 11773 246587
rect 12051 246309 29773 246587
rect 30051 246309 47773 246587
rect 48051 246309 65773 246587
rect 66051 246309 83773 246587
rect 84051 246309 101773 246587
rect 102051 246309 119773 246587
rect 120051 246309 137773 246587
rect 138051 246309 155773 246587
rect 156051 246309 173773 246587
rect 174051 246309 191773 246587
rect 192051 246309 209773 246587
rect 210051 246309 227773 246587
rect 228051 246309 245773 246587
rect 246051 246309 263773 246587
rect 264051 246309 281773 246587
rect 282051 246309 294111 246587
rect 294389 246309 294405 246587
rect -2443 246293 294405 246309
rect -1483 244727 293445 244743
rect -1483 244449 -1467 244727
rect -1189 244449 9913 244727
rect 10191 244449 27913 244727
rect 28191 244449 45913 244727
rect 46191 244449 63913 244727
rect 64191 244449 81913 244727
rect 82191 244449 99913 244727
rect 100191 244449 117913 244727
rect 118191 244449 135913 244727
rect 136191 244449 153913 244727
rect 154191 244449 171913 244727
rect 172191 244449 189913 244727
rect 190191 244449 207913 244727
rect 208191 244449 225913 244727
rect 226191 244449 243913 244727
rect 244191 244449 261913 244727
rect 262191 244449 279913 244727
rect 280191 244449 293151 244727
rect 293429 244449 293445 244727
rect -1483 244433 293445 244449
rect -4363 241307 296325 241323
rect -4363 241029 -3867 241307
rect -3589 241029 6493 241307
rect 6771 241029 24493 241307
rect 24771 241029 42493 241307
rect 42771 241029 60493 241307
rect 60771 241029 78493 241307
rect 78771 241029 96493 241307
rect 96771 241029 114493 241307
rect 114771 241029 132493 241307
rect 132771 241029 150493 241307
rect 150771 241029 168493 241307
rect 168771 241029 186493 241307
rect 186771 241029 204493 241307
rect 204771 241029 222493 241307
rect 222771 241029 240493 241307
rect 240771 241029 258493 241307
rect 258771 241029 276493 241307
rect 276771 241029 295551 241307
rect 295829 241029 296325 241307
rect -4363 241013 296325 241029
rect -3403 239447 295365 239463
rect -3403 239169 -2907 239447
rect -2629 239169 4633 239447
rect 4911 239169 22633 239447
rect 22911 239169 40633 239447
rect 40911 239169 58633 239447
rect 58911 239169 76633 239447
rect 76911 239169 94633 239447
rect 94911 239169 112633 239447
rect 112911 239169 130633 239447
rect 130911 239169 148633 239447
rect 148911 239169 166633 239447
rect 166911 239169 184633 239447
rect 184911 239169 202633 239447
rect 202911 239169 220633 239447
rect 220911 239169 238633 239447
rect 238911 239169 256633 239447
rect 256911 239169 274633 239447
rect 274911 239169 294591 239447
rect 294869 239169 295365 239447
rect -3403 239153 295365 239169
rect -2443 237587 294405 237603
rect -2443 237309 -1947 237587
rect -1669 237309 2773 237587
rect 3051 237309 20773 237587
rect 21051 237309 38773 237587
rect 39051 237309 56773 237587
rect 57051 237309 74773 237587
rect 75051 237309 92773 237587
rect 93051 237309 110773 237587
rect 111051 237309 128773 237587
rect 129051 237309 146773 237587
rect 147051 237309 164773 237587
rect 165051 237309 182773 237587
rect 183051 237309 200773 237587
rect 201051 237309 218773 237587
rect 219051 237309 236773 237587
rect 237051 237309 254773 237587
rect 255051 237309 272773 237587
rect 273051 237309 290773 237587
rect 291051 237309 293631 237587
rect 293909 237309 294405 237587
rect -2443 237293 294405 237309
rect -1483 235727 293445 235743
rect -1483 235449 -987 235727
rect -709 235449 913 235727
rect 1191 235449 18913 235727
rect 19191 235449 36913 235727
rect 37191 235449 54913 235727
rect 55191 235449 72913 235727
rect 73191 235449 90913 235727
rect 91191 235449 108913 235727
rect 109191 235449 126913 235727
rect 127191 235449 144913 235727
rect 145191 235449 162913 235727
rect 163191 235449 180913 235727
rect 181191 235449 198913 235727
rect 199191 235449 216913 235727
rect 217191 235449 234913 235727
rect 235191 235449 252913 235727
rect 253191 235449 270913 235727
rect 271191 235449 288913 235727
rect 289191 235449 292671 235727
rect 292949 235449 293445 235727
rect -1483 235433 293445 235449
rect -4363 232307 296325 232323
rect -4363 232029 -4347 232307
rect -4069 232029 15493 232307
rect 15771 232029 33493 232307
rect 33771 232029 51493 232307
rect 51771 232029 69493 232307
rect 69771 232029 87493 232307
rect 87771 232029 105493 232307
rect 105771 232029 123493 232307
rect 123771 232029 141493 232307
rect 141771 232029 159493 232307
rect 159771 232029 177493 232307
rect 177771 232029 195493 232307
rect 195771 232029 213493 232307
rect 213771 232029 231493 232307
rect 231771 232029 249493 232307
rect 249771 232029 267493 232307
rect 267771 232029 285493 232307
rect 285771 232029 296031 232307
rect 296309 232029 296325 232307
rect -4363 232013 296325 232029
rect -3403 230447 295365 230463
rect -3403 230169 -3387 230447
rect -3109 230169 13633 230447
rect 13911 230169 31633 230447
rect 31911 230169 49633 230447
rect 49911 230169 67633 230447
rect 67911 230169 85633 230447
rect 85911 230169 103633 230447
rect 103911 230169 121633 230447
rect 121911 230169 139633 230447
rect 139911 230169 157633 230447
rect 157911 230169 175633 230447
rect 175911 230169 193633 230447
rect 193911 230169 211633 230447
rect 211911 230169 229633 230447
rect 229911 230169 247633 230447
rect 247911 230169 265633 230447
rect 265911 230169 283633 230447
rect 283911 230169 295071 230447
rect 295349 230169 295365 230447
rect -3403 230153 295365 230169
rect -2443 228587 294405 228603
rect -2443 228309 -2427 228587
rect -2149 228309 11773 228587
rect 12051 228309 29773 228587
rect 30051 228309 47773 228587
rect 48051 228309 65773 228587
rect 66051 228309 83773 228587
rect 84051 228309 101773 228587
rect 102051 228309 119773 228587
rect 120051 228309 137773 228587
rect 138051 228309 155773 228587
rect 156051 228309 173773 228587
rect 174051 228309 191773 228587
rect 192051 228309 209773 228587
rect 210051 228309 227773 228587
rect 228051 228309 245773 228587
rect 246051 228309 263773 228587
rect 264051 228309 281773 228587
rect 282051 228309 294111 228587
rect 294389 228309 294405 228587
rect -2443 228293 294405 228309
rect -1483 226727 293445 226743
rect -1483 226449 -1467 226727
rect -1189 226449 9913 226727
rect 10191 226449 27913 226727
rect 28191 226449 45913 226727
rect 46191 226449 63913 226727
rect 64191 226449 81913 226727
rect 82191 226449 99913 226727
rect 100191 226449 117913 226727
rect 118191 226449 135913 226727
rect 136191 226449 153913 226727
rect 154191 226449 171913 226727
rect 172191 226449 189913 226727
rect 190191 226449 207913 226727
rect 208191 226449 225913 226727
rect 226191 226449 243913 226727
rect 244191 226449 261913 226727
rect 262191 226449 279913 226727
rect 280191 226449 293151 226727
rect 293429 226449 293445 226727
rect -1483 226433 293445 226449
rect -4363 223307 296325 223323
rect -4363 223029 -3867 223307
rect -3589 223029 6493 223307
rect 6771 223029 24493 223307
rect 24771 223029 42493 223307
rect 42771 223029 60493 223307
rect 60771 223029 78493 223307
rect 78771 223029 96493 223307
rect 96771 223029 114493 223307
rect 114771 223029 132493 223307
rect 132771 223029 150493 223307
rect 150771 223029 168493 223307
rect 168771 223029 186493 223307
rect 186771 223029 204493 223307
rect 204771 223029 222493 223307
rect 222771 223029 240493 223307
rect 240771 223029 258493 223307
rect 258771 223029 276493 223307
rect 276771 223029 295551 223307
rect 295829 223029 296325 223307
rect -4363 223013 296325 223029
rect -3403 221447 295365 221463
rect -3403 221169 -2907 221447
rect -2629 221169 4633 221447
rect 4911 221169 22633 221447
rect 22911 221169 40633 221447
rect 40911 221169 58633 221447
rect 58911 221169 76633 221447
rect 76911 221169 94633 221447
rect 94911 221169 112633 221447
rect 112911 221169 130633 221447
rect 130911 221169 148633 221447
rect 148911 221169 166633 221447
rect 166911 221169 184633 221447
rect 184911 221169 202633 221447
rect 202911 221169 220633 221447
rect 220911 221169 238633 221447
rect 238911 221169 256633 221447
rect 256911 221169 274633 221447
rect 274911 221169 294591 221447
rect 294869 221169 295365 221447
rect -3403 221153 295365 221169
rect -2443 219587 294405 219603
rect -2443 219309 -1947 219587
rect -1669 219309 2773 219587
rect 3051 219309 20773 219587
rect 21051 219309 38773 219587
rect 39051 219309 56773 219587
rect 57051 219309 74773 219587
rect 75051 219309 92773 219587
rect 93051 219309 110773 219587
rect 111051 219309 128773 219587
rect 129051 219309 146773 219587
rect 147051 219309 164773 219587
rect 165051 219309 182773 219587
rect 183051 219309 200773 219587
rect 201051 219309 218773 219587
rect 219051 219309 236773 219587
rect 237051 219309 254773 219587
rect 255051 219309 272773 219587
rect 273051 219309 290773 219587
rect 291051 219309 293631 219587
rect 293909 219309 294405 219587
rect -2443 219293 294405 219309
rect -1483 217727 293445 217743
rect -1483 217449 -987 217727
rect -709 217449 913 217727
rect 1191 217449 18913 217727
rect 19191 217449 36913 217727
rect 37191 217449 54913 217727
rect 55191 217449 72913 217727
rect 73191 217449 90913 217727
rect 91191 217449 108913 217727
rect 109191 217449 126913 217727
rect 127191 217449 144913 217727
rect 145191 217449 162913 217727
rect 163191 217449 180913 217727
rect 181191 217449 198913 217727
rect 199191 217449 216913 217727
rect 217191 217449 234913 217727
rect 235191 217449 252913 217727
rect 253191 217449 270913 217727
rect 271191 217449 288913 217727
rect 289191 217449 292671 217727
rect 292949 217449 293445 217727
rect -1483 217433 293445 217449
rect -4363 214307 296325 214323
rect -4363 214029 -4347 214307
rect -4069 214029 15493 214307
rect 15771 214029 33493 214307
rect 33771 214029 51493 214307
rect 51771 214029 69493 214307
rect 69771 214029 87493 214307
rect 87771 214029 105493 214307
rect 105771 214029 123493 214307
rect 123771 214029 141493 214307
rect 141771 214029 159493 214307
rect 159771 214029 177493 214307
rect 177771 214029 195493 214307
rect 195771 214029 213493 214307
rect 213771 214029 231493 214307
rect 231771 214029 249493 214307
rect 249771 214029 267493 214307
rect 267771 214029 285493 214307
rect 285771 214029 296031 214307
rect 296309 214029 296325 214307
rect -4363 214013 296325 214029
rect -3403 212447 295365 212463
rect -3403 212169 -3387 212447
rect -3109 212169 13633 212447
rect 13911 212169 31633 212447
rect 31911 212169 49633 212447
rect 49911 212169 67633 212447
rect 67911 212169 85633 212447
rect 85911 212169 103633 212447
rect 103911 212169 121633 212447
rect 121911 212169 139633 212447
rect 139911 212169 157633 212447
rect 157911 212169 175633 212447
rect 175911 212169 193633 212447
rect 193911 212169 211633 212447
rect 211911 212169 229633 212447
rect 229911 212169 247633 212447
rect 247911 212169 265633 212447
rect 265911 212169 283633 212447
rect 283911 212169 295071 212447
rect 295349 212169 295365 212447
rect -3403 212153 295365 212169
rect -2443 210587 294405 210603
rect -2443 210309 -2427 210587
rect -2149 210309 11773 210587
rect 12051 210309 29773 210587
rect 30051 210309 47773 210587
rect 48051 210309 65773 210587
rect 66051 210309 83773 210587
rect 84051 210309 101773 210587
rect 102051 210309 119773 210587
rect 120051 210309 137773 210587
rect 138051 210309 155773 210587
rect 156051 210309 173773 210587
rect 174051 210309 191773 210587
rect 192051 210309 209773 210587
rect 210051 210309 227773 210587
rect 228051 210309 245773 210587
rect 246051 210309 263773 210587
rect 264051 210309 281773 210587
rect 282051 210309 294111 210587
rect 294389 210309 294405 210587
rect -2443 210293 294405 210309
rect -1483 208727 293445 208743
rect -1483 208449 -1467 208727
rect -1189 208449 9913 208727
rect 10191 208449 27913 208727
rect 28191 208449 45913 208727
rect 46191 208449 63913 208727
rect 64191 208449 81913 208727
rect 82191 208449 99913 208727
rect 100191 208449 117913 208727
rect 118191 208449 135913 208727
rect 136191 208449 153913 208727
rect 154191 208449 171913 208727
rect 172191 208449 189913 208727
rect 190191 208449 207913 208727
rect 208191 208449 225913 208727
rect 226191 208449 243913 208727
rect 244191 208449 261913 208727
rect 262191 208449 279913 208727
rect 280191 208449 293151 208727
rect 293429 208449 293445 208727
rect -1483 208433 293445 208449
rect -4363 205307 296325 205323
rect -4363 205029 -3867 205307
rect -3589 205029 6493 205307
rect 6771 205029 24493 205307
rect 24771 205029 42493 205307
rect 42771 205029 60493 205307
rect 60771 205029 78493 205307
rect 78771 205029 96493 205307
rect 96771 205029 114493 205307
rect 114771 205029 132493 205307
rect 132771 205029 150493 205307
rect 150771 205029 168493 205307
rect 168771 205029 186493 205307
rect 186771 205029 204493 205307
rect 204771 205029 222493 205307
rect 222771 205029 240493 205307
rect 240771 205029 258493 205307
rect 258771 205029 276493 205307
rect 276771 205029 295551 205307
rect 295829 205029 296325 205307
rect -4363 205013 296325 205029
rect -3403 203447 295365 203463
rect -3403 203169 -2907 203447
rect -2629 203169 4633 203447
rect 4911 203169 22633 203447
rect 22911 203169 40633 203447
rect 40911 203169 58633 203447
rect 58911 203169 76633 203447
rect 76911 203169 94633 203447
rect 94911 203169 112633 203447
rect 112911 203169 130633 203447
rect 130911 203169 148633 203447
rect 148911 203169 166633 203447
rect 166911 203169 184633 203447
rect 184911 203169 202633 203447
rect 202911 203169 220633 203447
rect 220911 203169 238633 203447
rect 238911 203169 256633 203447
rect 256911 203169 274633 203447
rect 274911 203169 294591 203447
rect 294869 203169 295365 203447
rect -3403 203153 295365 203169
rect -2443 201587 294405 201603
rect -2443 201309 -1947 201587
rect -1669 201309 2773 201587
rect 3051 201309 20773 201587
rect 21051 201309 38773 201587
rect 39051 201309 56773 201587
rect 57051 201309 74773 201587
rect 75051 201309 92773 201587
rect 93051 201309 110773 201587
rect 111051 201309 128773 201587
rect 129051 201309 146773 201587
rect 147051 201309 164773 201587
rect 165051 201309 182773 201587
rect 183051 201309 200773 201587
rect 201051 201309 218773 201587
rect 219051 201309 236773 201587
rect 237051 201309 254773 201587
rect 255051 201309 272773 201587
rect 273051 201309 290773 201587
rect 291051 201309 293631 201587
rect 293909 201309 294405 201587
rect -2443 201293 294405 201309
rect -1483 199727 293445 199743
rect -1483 199449 -987 199727
rect -709 199449 913 199727
rect 1191 199449 18913 199727
rect 19191 199449 36913 199727
rect 37191 199449 54913 199727
rect 55191 199449 72913 199727
rect 73191 199449 90913 199727
rect 91191 199449 108913 199727
rect 109191 199449 126913 199727
rect 127191 199449 144913 199727
rect 145191 199449 162913 199727
rect 163191 199449 180913 199727
rect 181191 199449 198913 199727
rect 199191 199449 216913 199727
rect 217191 199449 234913 199727
rect 235191 199449 252913 199727
rect 253191 199449 270913 199727
rect 271191 199449 288913 199727
rect 289191 199449 292671 199727
rect 292949 199449 293445 199727
rect -1483 199433 293445 199449
rect -4363 196307 296325 196323
rect -4363 196029 -4347 196307
rect -4069 196029 15493 196307
rect 15771 196029 33493 196307
rect 33771 196029 51493 196307
rect 51771 196029 69493 196307
rect 69771 196029 87493 196307
rect 87771 196029 105493 196307
rect 105771 196029 123493 196307
rect 123771 196029 141493 196307
rect 141771 196029 159493 196307
rect 159771 196029 177493 196307
rect 177771 196029 195493 196307
rect 195771 196029 213493 196307
rect 213771 196029 231493 196307
rect 231771 196029 249493 196307
rect 249771 196029 267493 196307
rect 267771 196029 285493 196307
rect 285771 196029 296031 196307
rect 296309 196029 296325 196307
rect -4363 196013 296325 196029
rect -3403 194447 295365 194463
rect -3403 194169 -3387 194447
rect -3109 194169 13633 194447
rect 13911 194169 31633 194447
rect 31911 194169 49633 194447
rect 49911 194169 67633 194447
rect 67911 194169 85633 194447
rect 85911 194169 103633 194447
rect 103911 194169 121633 194447
rect 121911 194169 139633 194447
rect 139911 194169 157633 194447
rect 157911 194169 175633 194447
rect 175911 194169 193633 194447
rect 193911 194169 211633 194447
rect 211911 194169 229633 194447
rect 229911 194169 247633 194447
rect 247911 194169 265633 194447
rect 265911 194169 283633 194447
rect 283911 194169 295071 194447
rect 295349 194169 295365 194447
rect -3403 194153 295365 194169
rect -2443 192587 294405 192603
rect -2443 192309 -2427 192587
rect -2149 192309 11773 192587
rect 12051 192309 29773 192587
rect 30051 192309 47773 192587
rect 48051 192309 65773 192587
rect 66051 192309 83773 192587
rect 84051 192309 101773 192587
rect 102051 192309 119773 192587
rect 120051 192309 137773 192587
rect 138051 192309 155773 192587
rect 156051 192309 173773 192587
rect 174051 192309 191773 192587
rect 192051 192309 209773 192587
rect 210051 192309 227773 192587
rect 228051 192309 245773 192587
rect 246051 192309 263773 192587
rect 264051 192309 281773 192587
rect 282051 192309 294111 192587
rect 294389 192309 294405 192587
rect -2443 192293 294405 192309
rect -1483 190727 293445 190743
rect -1483 190449 -1467 190727
rect -1189 190449 9913 190727
rect 10191 190449 27913 190727
rect 28191 190449 45913 190727
rect 46191 190449 63913 190727
rect 64191 190449 81913 190727
rect 82191 190449 99913 190727
rect 100191 190449 117913 190727
rect 118191 190449 135913 190727
rect 136191 190449 153913 190727
rect 154191 190449 171913 190727
rect 172191 190449 189913 190727
rect 190191 190449 207913 190727
rect 208191 190449 225913 190727
rect 226191 190449 243913 190727
rect 244191 190449 261913 190727
rect 262191 190449 279913 190727
rect 280191 190449 293151 190727
rect 293429 190449 293445 190727
rect -1483 190433 293445 190449
rect -4363 187307 296325 187323
rect -4363 187029 -3867 187307
rect -3589 187029 6493 187307
rect 6771 187029 24493 187307
rect 24771 187029 42493 187307
rect 42771 187029 60493 187307
rect 60771 187029 78493 187307
rect 78771 187029 96493 187307
rect 96771 187029 114493 187307
rect 114771 187029 132493 187307
rect 132771 187029 150493 187307
rect 150771 187029 168493 187307
rect 168771 187029 186493 187307
rect 186771 187029 204493 187307
rect 204771 187029 222493 187307
rect 222771 187029 240493 187307
rect 240771 187029 258493 187307
rect 258771 187029 276493 187307
rect 276771 187029 295551 187307
rect 295829 187029 296325 187307
rect -4363 187013 296325 187029
rect -3403 185447 295365 185463
rect -3403 185169 -2907 185447
rect -2629 185169 4633 185447
rect 4911 185169 22633 185447
rect 22911 185169 40633 185447
rect 40911 185169 58633 185447
rect 58911 185169 76633 185447
rect 76911 185169 94633 185447
rect 94911 185169 112633 185447
rect 112911 185169 130633 185447
rect 130911 185169 148633 185447
rect 148911 185169 166633 185447
rect 166911 185169 184633 185447
rect 184911 185169 202633 185447
rect 202911 185169 220633 185447
rect 220911 185169 238633 185447
rect 238911 185169 256633 185447
rect 256911 185169 274633 185447
rect 274911 185169 294591 185447
rect 294869 185169 295365 185447
rect -3403 185153 295365 185169
rect -2443 183587 294405 183603
rect -2443 183309 -1947 183587
rect -1669 183309 2773 183587
rect 3051 183309 20773 183587
rect 21051 183309 38773 183587
rect 39051 183309 56773 183587
rect 57051 183309 74773 183587
rect 75051 183309 92773 183587
rect 93051 183309 110773 183587
rect 111051 183309 128773 183587
rect 129051 183309 146773 183587
rect 147051 183309 164773 183587
rect 165051 183309 182773 183587
rect 183051 183309 200773 183587
rect 201051 183309 218773 183587
rect 219051 183309 236773 183587
rect 237051 183309 254773 183587
rect 255051 183309 272773 183587
rect 273051 183309 290773 183587
rect 291051 183309 293631 183587
rect 293909 183309 294405 183587
rect -2443 183293 294405 183309
rect -1483 181727 293445 181743
rect -1483 181449 -987 181727
rect -709 181449 913 181727
rect 1191 181449 18913 181727
rect 19191 181449 36913 181727
rect 37191 181449 54913 181727
rect 55191 181449 72913 181727
rect 73191 181449 90913 181727
rect 91191 181449 108913 181727
rect 109191 181449 126913 181727
rect 127191 181449 144913 181727
rect 145191 181449 162913 181727
rect 163191 181449 180913 181727
rect 181191 181449 198913 181727
rect 199191 181449 216913 181727
rect 217191 181449 234913 181727
rect 235191 181449 252913 181727
rect 253191 181449 270913 181727
rect 271191 181449 288913 181727
rect 289191 181449 292671 181727
rect 292949 181449 293445 181727
rect -1483 181433 293445 181449
rect -4363 178307 296325 178323
rect -4363 178029 -4347 178307
rect -4069 178029 15493 178307
rect 15771 178029 33493 178307
rect 33771 178029 51493 178307
rect 51771 178029 69493 178307
rect 69771 178029 87493 178307
rect 87771 178029 105493 178307
rect 105771 178029 123493 178307
rect 123771 178029 141493 178307
rect 141771 178029 159493 178307
rect 159771 178029 177493 178307
rect 177771 178029 195493 178307
rect 195771 178029 213493 178307
rect 213771 178029 231493 178307
rect 231771 178029 249493 178307
rect 249771 178029 267493 178307
rect 267771 178029 285493 178307
rect 285771 178029 296031 178307
rect 296309 178029 296325 178307
rect -4363 178013 296325 178029
rect -3403 176447 295365 176463
rect -3403 176169 -3387 176447
rect -3109 176169 13633 176447
rect 13911 176169 31633 176447
rect 31911 176169 49633 176447
rect 49911 176169 67633 176447
rect 67911 176169 85633 176447
rect 85911 176169 103633 176447
rect 103911 176169 121633 176447
rect 121911 176169 139633 176447
rect 139911 176169 157633 176447
rect 157911 176169 175633 176447
rect 175911 176169 193633 176447
rect 193911 176169 211633 176447
rect 211911 176169 229633 176447
rect 229911 176169 247633 176447
rect 247911 176169 265633 176447
rect 265911 176169 283633 176447
rect 283911 176169 295071 176447
rect 295349 176169 295365 176447
rect -3403 176153 295365 176169
rect -2443 174587 294405 174603
rect -2443 174309 -2427 174587
rect -2149 174309 11773 174587
rect 12051 174309 29773 174587
rect 30051 174309 47773 174587
rect 48051 174309 65773 174587
rect 66051 174309 83773 174587
rect 84051 174309 101773 174587
rect 102051 174309 119773 174587
rect 120051 174309 137773 174587
rect 138051 174309 155773 174587
rect 156051 174309 173773 174587
rect 174051 174309 191773 174587
rect 192051 174309 209773 174587
rect 210051 174309 227773 174587
rect 228051 174309 245773 174587
rect 246051 174309 263773 174587
rect 264051 174309 281773 174587
rect 282051 174309 294111 174587
rect 294389 174309 294405 174587
rect -2443 174293 294405 174309
rect -1483 172727 293445 172743
rect -1483 172449 -1467 172727
rect -1189 172449 9913 172727
rect 10191 172449 27913 172727
rect 28191 172449 45913 172727
rect 46191 172449 63913 172727
rect 64191 172449 81913 172727
rect 82191 172449 99913 172727
rect 100191 172449 117913 172727
rect 118191 172449 135913 172727
rect 136191 172449 153913 172727
rect 154191 172449 171913 172727
rect 172191 172449 189913 172727
rect 190191 172449 207913 172727
rect 208191 172449 225913 172727
rect 226191 172449 243913 172727
rect 244191 172449 261913 172727
rect 262191 172449 279913 172727
rect 280191 172449 293151 172727
rect 293429 172449 293445 172727
rect -1483 172433 293445 172449
rect -4363 169307 296325 169323
rect -4363 169029 -3867 169307
rect -3589 169029 6493 169307
rect 6771 169029 24493 169307
rect 24771 169029 42493 169307
rect 42771 169029 60493 169307
rect 60771 169029 78493 169307
rect 78771 169029 96493 169307
rect 96771 169029 114493 169307
rect 114771 169029 132493 169307
rect 132771 169029 150493 169307
rect 150771 169029 168493 169307
rect 168771 169029 186493 169307
rect 186771 169029 204493 169307
rect 204771 169029 222493 169307
rect 222771 169029 240493 169307
rect 240771 169029 258493 169307
rect 258771 169029 276493 169307
rect 276771 169029 295551 169307
rect 295829 169029 296325 169307
rect -4363 169013 296325 169029
rect -3403 167447 295365 167463
rect -3403 167169 -2907 167447
rect -2629 167169 4633 167447
rect 4911 167169 22633 167447
rect 22911 167169 40633 167447
rect 40911 167169 58633 167447
rect 58911 167169 76633 167447
rect 76911 167169 94633 167447
rect 94911 167169 112633 167447
rect 112911 167169 130633 167447
rect 130911 167169 148633 167447
rect 148911 167169 166633 167447
rect 166911 167169 184633 167447
rect 184911 167169 202633 167447
rect 202911 167169 220633 167447
rect 220911 167169 238633 167447
rect 238911 167169 256633 167447
rect 256911 167169 274633 167447
rect 274911 167169 294591 167447
rect 294869 167169 295365 167447
rect -3403 167153 295365 167169
rect -2443 165587 294405 165603
rect -2443 165309 -1947 165587
rect -1669 165309 2773 165587
rect 3051 165309 20773 165587
rect 21051 165309 38773 165587
rect 39051 165309 56773 165587
rect 57051 165309 74773 165587
rect 75051 165309 92773 165587
rect 93051 165309 110773 165587
rect 111051 165309 128773 165587
rect 129051 165309 146773 165587
rect 147051 165309 164773 165587
rect 165051 165309 182773 165587
rect 183051 165309 200773 165587
rect 201051 165309 218773 165587
rect 219051 165309 236773 165587
rect 237051 165309 254773 165587
rect 255051 165309 272773 165587
rect 273051 165309 290773 165587
rect 291051 165309 293631 165587
rect 293909 165309 294405 165587
rect -2443 165293 294405 165309
rect -1483 163727 293445 163743
rect -1483 163449 -987 163727
rect -709 163449 913 163727
rect 1191 163449 18913 163727
rect 19191 163449 36913 163727
rect 37191 163449 54913 163727
rect 55191 163449 72913 163727
rect 73191 163449 90913 163727
rect 91191 163449 108913 163727
rect 109191 163449 126913 163727
rect 127191 163449 144913 163727
rect 145191 163449 162913 163727
rect 163191 163449 180913 163727
rect 181191 163449 198913 163727
rect 199191 163449 216913 163727
rect 217191 163449 234913 163727
rect 235191 163449 252913 163727
rect 253191 163449 270913 163727
rect 271191 163449 288913 163727
rect 289191 163449 292671 163727
rect 292949 163449 293445 163727
rect -1483 163433 293445 163449
rect -4363 160307 296325 160323
rect -4363 160029 -4347 160307
rect -4069 160029 15493 160307
rect 15771 160029 33493 160307
rect 33771 160029 51493 160307
rect 51771 160029 69493 160307
rect 69771 160029 87493 160307
rect 87771 160029 105493 160307
rect 105771 160029 123493 160307
rect 123771 160029 141493 160307
rect 141771 160029 159493 160307
rect 159771 160029 177493 160307
rect 177771 160029 195493 160307
rect 195771 160029 213493 160307
rect 213771 160029 231493 160307
rect 231771 160029 249493 160307
rect 249771 160029 267493 160307
rect 267771 160029 285493 160307
rect 285771 160029 296031 160307
rect 296309 160029 296325 160307
rect -4363 160013 296325 160029
rect -3403 158447 295365 158463
rect -3403 158169 -3387 158447
rect -3109 158169 13633 158447
rect 13911 158169 31633 158447
rect 31911 158169 49633 158447
rect 49911 158169 67633 158447
rect 67911 158169 85633 158447
rect 85911 158169 103633 158447
rect 103911 158169 121633 158447
rect 121911 158169 139633 158447
rect 139911 158169 157633 158447
rect 157911 158169 175633 158447
rect 175911 158169 193633 158447
rect 193911 158169 211633 158447
rect 211911 158169 229633 158447
rect 229911 158169 247633 158447
rect 247911 158169 265633 158447
rect 265911 158169 283633 158447
rect 283911 158169 295071 158447
rect 295349 158169 295365 158447
rect -3403 158153 295365 158169
rect -2443 156587 294405 156603
rect -2443 156309 -2427 156587
rect -2149 156309 11773 156587
rect 12051 156309 29773 156587
rect 30051 156309 47773 156587
rect 48051 156309 65773 156587
rect 66051 156309 83773 156587
rect 84051 156309 101773 156587
rect 102051 156309 119773 156587
rect 120051 156309 137773 156587
rect 138051 156309 155773 156587
rect 156051 156309 173773 156587
rect 174051 156309 191773 156587
rect 192051 156309 209773 156587
rect 210051 156309 227773 156587
rect 228051 156309 245773 156587
rect 246051 156309 263773 156587
rect 264051 156309 281773 156587
rect 282051 156309 294111 156587
rect 294389 156309 294405 156587
rect -2443 156293 294405 156309
rect -1483 154727 293445 154743
rect -1483 154449 -1467 154727
rect -1189 154449 9913 154727
rect 10191 154449 27913 154727
rect 28191 154449 45913 154727
rect 46191 154449 63913 154727
rect 64191 154449 81913 154727
rect 82191 154449 99913 154727
rect 100191 154449 117913 154727
rect 118191 154449 135913 154727
rect 136191 154449 153913 154727
rect 154191 154449 171913 154727
rect 172191 154449 189913 154727
rect 190191 154449 207913 154727
rect 208191 154449 225913 154727
rect 226191 154449 243913 154727
rect 244191 154449 261913 154727
rect 262191 154449 279913 154727
rect 280191 154449 293151 154727
rect 293429 154449 293445 154727
rect -1483 154433 293445 154449
rect -4363 151307 296325 151323
rect -4363 151029 -3867 151307
rect -3589 151029 6493 151307
rect 6771 151029 24493 151307
rect 24771 151029 42493 151307
rect 42771 151029 60493 151307
rect 60771 151029 78493 151307
rect 78771 151029 96493 151307
rect 96771 151029 114493 151307
rect 114771 151029 132493 151307
rect 132771 151029 150493 151307
rect 150771 151029 168493 151307
rect 168771 151029 186493 151307
rect 186771 151029 204493 151307
rect 204771 151029 222493 151307
rect 222771 151029 240493 151307
rect 240771 151029 258493 151307
rect 258771 151029 276493 151307
rect 276771 151029 295551 151307
rect 295829 151029 296325 151307
rect -4363 151013 296325 151029
rect -3403 149447 295365 149463
rect -3403 149169 -2907 149447
rect -2629 149169 4633 149447
rect 4911 149169 22633 149447
rect 22911 149169 40633 149447
rect 40911 149169 58633 149447
rect 58911 149169 76633 149447
rect 76911 149169 94633 149447
rect 94911 149169 112633 149447
rect 112911 149169 130633 149447
rect 130911 149169 148633 149447
rect 148911 149169 166633 149447
rect 166911 149169 184633 149447
rect 184911 149169 202633 149447
rect 202911 149169 220633 149447
rect 220911 149169 238633 149447
rect 238911 149169 256633 149447
rect 256911 149169 274633 149447
rect 274911 149169 294591 149447
rect 294869 149169 295365 149447
rect -3403 149153 295365 149169
rect -2443 147587 294405 147603
rect -2443 147309 -1947 147587
rect -1669 147309 2773 147587
rect 3051 147309 20773 147587
rect 21051 147309 38773 147587
rect 39051 147309 56773 147587
rect 57051 147309 74773 147587
rect 75051 147309 92773 147587
rect 93051 147309 110773 147587
rect 111051 147309 128773 147587
rect 129051 147309 146773 147587
rect 147051 147309 164773 147587
rect 165051 147309 182773 147587
rect 183051 147309 200773 147587
rect 201051 147309 218773 147587
rect 219051 147309 236773 147587
rect 237051 147309 254773 147587
rect 255051 147309 272773 147587
rect 273051 147309 290773 147587
rect 291051 147309 293631 147587
rect 293909 147309 294405 147587
rect -2443 147293 294405 147309
rect -1483 145727 293445 145743
rect -1483 145449 -987 145727
rect -709 145449 913 145727
rect 1191 145449 18913 145727
rect 19191 145449 36913 145727
rect 37191 145449 54913 145727
rect 55191 145449 72913 145727
rect 73191 145449 90913 145727
rect 91191 145449 108913 145727
rect 109191 145449 126913 145727
rect 127191 145449 144913 145727
rect 145191 145449 162913 145727
rect 163191 145449 180913 145727
rect 181191 145449 198913 145727
rect 199191 145449 216913 145727
rect 217191 145449 234913 145727
rect 235191 145449 252913 145727
rect 253191 145449 270913 145727
rect 271191 145449 288913 145727
rect 289191 145449 292671 145727
rect 292949 145449 293445 145727
rect -1483 145433 293445 145449
rect -4363 142307 296325 142323
rect -4363 142029 -4347 142307
rect -4069 142029 15493 142307
rect 15771 142029 33493 142307
rect 33771 142029 51493 142307
rect 51771 142029 69493 142307
rect 69771 142029 87493 142307
rect 87771 142029 105493 142307
rect 105771 142029 123493 142307
rect 123771 142029 141493 142307
rect 141771 142029 159493 142307
rect 159771 142029 177493 142307
rect 177771 142029 195493 142307
rect 195771 142029 213493 142307
rect 213771 142029 231493 142307
rect 231771 142029 249493 142307
rect 249771 142029 267493 142307
rect 267771 142029 285493 142307
rect 285771 142029 296031 142307
rect 296309 142029 296325 142307
rect -4363 142013 296325 142029
rect -3403 140447 295365 140463
rect -3403 140169 -3387 140447
rect -3109 140169 13633 140447
rect 13911 140169 31633 140447
rect 31911 140169 49633 140447
rect 49911 140169 67633 140447
rect 67911 140169 85633 140447
rect 85911 140169 103633 140447
rect 103911 140169 121633 140447
rect 121911 140169 139633 140447
rect 139911 140169 157633 140447
rect 157911 140169 175633 140447
rect 175911 140169 193633 140447
rect 193911 140169 211633 140447
rect 211911 140169 229633 140447
rect 229911 140169 247633 140447
rect 247911 140169 265633 140447
rect 265911 140169 283633 140447
rect 283911 140169 295071 140447
rect 295349 140169 295365 140447
rect -3403 140153 295365 140169
rect -2443 138587 294405 138603
rect -2443 138309 -2427 138587
rect -2149 138309 11773 138587
rect 12051 138309 29773 138587
rect 30051 138309 47773 138587
rect 48051 138309 65773 138587
rect 66051 138309 83773 138587
rect 84051 138309 101773 138587
rect 102051 138309 119773 138587
rect 120051 138309 137773 138587
rect 138051 138309 155773 138587
rect 156051 138309 173773 138587
rect 174051 138309 191773 138587
rect 192051 138309 209773 138587
rect 210051 138309 227773 138587
rect 228051 138309 245773 138587
rect 246051 138309 263773 138587
rect 264051 138309 281773 138587
rect 282051 138309 294111 138587
rect 294389 138309 294405 138587
rect -2443 138293 294405 138309
rect -1483 136727 293445 136743
rect -1483 136449 -1467 136727
rect -1189 136449 9913 136727
rect 10191 136449 27913 136727
rect 28191 136449 45913 136727
rect 46191 136449 63913 136727
rect 64191 136449 81913 136727
rect 82191 136449 99913 136727
rect 100191 136449 117913 136727
rect 118191 136449 135913 136727
rect 136191 136449 153913 136727
rect 154191 136449 171913 136727
rect 172191 136449 189913 136727
rect 190191 136449 207913 136727
rect 208191 136449 225913 136727
rect 226191 136449 243913 136727
rect 244191 136449 261913 136727
rect 262191 136449 279913 136727
rect 280191 136449 293151 136727
rect 293429 136449 293445 136727
rect -1483 136433 293445 136449
rect -4363 133307 296325 133323
rect -4363 133029 -3867 133307
rect -3589 133029 6493 133307
rect 6771 133029 24493 133307
rect 24771 133029 42493 133307
rect 42771 133029 60493 133307
rect 60771 133029 78493 133307
rect 78771 133029 96493 133307
rect 96771 133029 114493 133307
rect 114771 133029 132493 133307
rect 132771 133029 150493 133307
rect 150771 133029 168493 133307
rect 168771 133029 186493 133307
rect 186771 133029 204493 133307
rect 204771 133029 222493 133307
rect 222771 133029 240493 133307
rect 240771 133029 258493 133307
rect 258771 133029 276493 133307
rect 276771 133029 295551 133307
rect 295829 133029 296325 133307
rect -4363 133013 296325 133029
rect -3403 131447 295365 131463
rect -3403 131169 -2907 131447
rect -2629 131169 4633 131447
rect 4911 131169 22633 131447
rect 22911 131169 40633 131447
rect 40911 131169 58633 131447
rect 58911 131169 76633 131447
rect 76911 131169 94633 131447
rect 94911 131169 112633 131447
rect 112911 131169 130633 131447
rect 130911 131169 148633 131447
rect 148911 131169 166633 131447
rect 166911 131169 184633 131447
rect 184911 131169 202633 131447
rect 202911 131169 220633 131447
rect 220911 131169 238633 131447
rect 238911 131169 256633 131447
rect 256911 131169 274633 131447
rect 274911 131169 294591 131447
rect 294869 131169 295365 131447
rect -3403 131153 295365 131169
rect -2443 129587 294405 129603
rect -2443 129309 -1947 129587
rect -1669 129309 2773 129587
rect 3051 129309 20773 129587
rect 21051 129309 38773 129587
rect 39051 129309 56773 129587
rect 57051 129309 74773 129587
rect 75051 129309 92773 129587
rect 93051 129309 110773 129587
rect 111051 129309 128773 129587
rect 129051 129309 146773 129587
rect 147051 129309 164773 129587
rect 165051 129309 182773 129587
rect 183051 129309 200773 129587
rect 201051 129309 218773 129587
rect 219051 129309 236773 129587
rect 237051 129309 254773 129587
rect 255051 129309 272773 129587
rect 273051 129309 290773 129587
rect 291051 129309 293631 129587
rect 293909 129309 294405 129587
rect -2443 129293 294405 129309
rect -1483 127727 293445 127743
rect -1483 127449 -987 127727
rect -709 127449 913 127727
rect 1191 127449 18913 127727
rect 19191 127449 36913 127727
rect 37191 127449 54913 127727
rect 55191 127449 72913 127727
rect 73191 127449 90913 127727
rect 91191 127449 108913 127727
rect 109191 127449 126913 127727
rect 127191 127449 144913 127727
rect 145191 127449 162913 127727
rect 163191 127449 180913 127727
rect 181191 127449 198913 127727
rect 199191 127449 216913 127727
rect 217191 127449 234913 127727
rect 235191 127449 252913 127727
rect 253191 127449 270913 127727
rect 271191 127449 288913 127727
rect 289191 127449 292671 127727
rect 292949 127449 293445 127727
rect -1483 127433 293445 127449
rect -4363 124307 296325 124323
rect -4363 124029 -4347 124307
rect -4069 124029 15493 124307
rect 15771 124029 33493 124307
rect 33771 124029 51493 124307
rect 51771 124029 69493 124307
rect 69771 124029 87493 124307
rect 87771 124029 105493 124307
rect 105771 124029 123493 124307
rect 123771 124029 141493 124307
rect 141771 124029 159493 124307
rect 159771 124029 177493 124307
rect 177771 124029 195493 124307
rect 195771 124029 213493 124307
rect 213771 124029 231493 124307
rect 231771 124029 249493 124307
rect 249771 124029 267493 124307
rect 267771 124029 285493 124307
rect 285771 124029 296031 124307
rect 296309 124029 296325 124307
rect -4363 124013 296325 124029
rect -3403 122447 295365 122463
rect -3403 122169 -3387 122447
rect -3109 122169 13633 122447
rect 13911 122169 31633 122447
rect 31911 122169 49633 122447
rect 49911 122169 67633 122447
rect 67911 122169 85633 122447
rect 85911 122169 103633 122447
rect 103911 122169 121633 122447
rect 121911 122169 139633 122447
rect 139911 122169 157633 122447
rect 157911 122169 175633 122447
rect 175911 122169 193633 122447
rect 193911 122169 211633 122447
rect 211911 122169 229633 122447
rect 229911 122169 247633 122447
rect 247911 122169 265633 122447
rect 265911 122169 283633 122447
rect 283911 122169 295071 122447
rect 295349 122169 295365 122447
rect -3403 122153 295365 122169
rect -2443 120587 294405 120603
rect -2443 120309 -2427 120587
rect -2149 120309 11773 120587
rect 12051 120309 29773 120587
rect 30051 120309 47773 120587
rect 48051 120309 65773 120587
rect 66051 120309 83773 120587
rect 84051 120309 101773 120587
rect 102051 120309 119773 120587
rect 120051 120309 137773 120587
rect 138051 120309 155773 120587
rect 156051 120309 173773 120587
rect 174051 120309 191773 120587
rect 192051 120309 209773 120587
rect 210051 120309 227773 120587
rect 228051 120309 245773 120587
rect 246051 120309 263773 120587
rect 264051 120309 281773 120587
rect 282051 120309 294111 120587
rect 294389 120309 294405 120587
rect -2443 120293 294405 120309
rect -1483 118727 293445 118743
rect -1483 118449 -1467 118727
rect -1189 118449 9913 118727
rect 10191 118449 27913 118727
rect 28191 118449 45913 118727
rect 46191 118449 63913 118727
rect 64191 118449 81913 118727
rect 82191 118449 99913 118727
rect 100191 118449 117913 118727
rect 118191 118449 135913 118727
rect 136191 118449 153913 118727
rect 154191 118449 171913 118727
rect 172191 118449 189913 118727
rect 190191 118449 207913 118727
rect 208191 118449 225913 118727
rect 226191 118449 243913 118727
rect 244191 118449 261913 118727
rect 262191 118449 279913 118727
rect 280191 118449 293151 118727
rect 293429 118449 293445 118727
rect -1483 118433 293445 118449
rect -4363 115307 296325 115323
rect -4363 115029 -3867 115307
rect -3589 115029 6493 115307
rect 6771 115029 24493 115307
rect 24771 115029 42493 115307
rect 42771 115029 60493 115307
rect 60771 115029 78493 115307
rect 78771 115029 96493 115307
rect 96771 115029 114493 115307
rect 114771 115029 132493 115307
rect 132771 115029 150493 115307
rect 150771 115029 168493 115307
rect 168771 115029 186493 115307
rect 186771 115029 204493 115307
rect 204771 115029 222493 115307
rect 222771 115029 240493 115307
rect 240771 115029 258493 115307
rect 258771 115029 276493 115307
rect 276771 115029 295551 115307
rect 295829 115029 296325 115307
rect -4363 115013 296325 115029
rect -3403 113447 295365 113463
rect -3403 113169 -2907 113447
rect -2629 113169 4633 113447
rect 4911 113169 22633 113447
rect 22911 113169 40633 113447
rect 40911 113169 58633 113447
rect 58911 113169 76633 113447
rect 76911 113169 94633 113447
rect 94911 113169 112633 113447
rect 112911 113169 130633 113447
rect 130911 113169 148633 113447
rect 148911 113169 166633 113447
rect 166911 113169 184633 113447
rect 184911 113169 202633 113447
rect 202911 113169 220633 113447
rect 220911 113169 238633 113447
rect 238911 113169 256633 113447
rect 256911 113169 274633 113447
rect 274911 113169 294591 113447
rect 294869 113169 295365 113447
rect -3403 113153 295365 113169
rect -2443 111587 294405 111603
rect -2443 111309 -1947 111587
rect -1669 111309 2773 111587
rect 3051 111309 20773 111587
rect 21051 111309 38773 111587
rect 39051 111309 56773 111587
rect 57051 111309 74773 111587
rect 75051 111309 92773 111587
rect 93051 111309 110773 111587
rect 111051 111309 128773 111587
rect 129051 111309 146773 111587
rect 147051 111309 164773 111587
rect 165051 111309 182773 111587
rect 183051 111309 200773 111587
rect 201051 111309 218773 111587
rect 219051 111309 236773 111587
rect 237051 111309 254773 111587
rect 255051 111309 272773 111587
rect 273051 111309 290773 111587
rect 291051 111309 293631 111587
rect 293909 111309 294405 111587
rect -2443 111293 294405 111309
rect -1483 109727 293445 109743
rect -1483 109449 -987 109727
rect -709 109449 913 109727
rect 1191 109449 18913 109727
rect 19191 109449 36913 109727
rect 37191 109449 54913 109727
rect 55191 109449 72913 109727
rect 73191 109449 90913 109727
rect 91191 109449 108913 109727
rect 109191 109449 126913 109727
rect 127191 109449 144913 109727
rect 145191 109449 162913 109727
rect 163191 109449 180913 109727
rect 181191 109449 198913 109727
rect 199191 109449 216913 109727
rect 217191 109449 234913 109727
rect 235191 109449 252913 109727
rect 253191 109449 270913 109727
rect 271191 109449 288913 109727
rect 289191 109449 292671 109727
rect 292949 109449 293445 109727
rect -1483 109433 293445 109449
rect -4363 106307 296325 106323
rect -4363 106029 -4347 106307
rect -4069 106029 15493 106307
rect 15771 106029 33493 106307
rect 33771 106029 51493 106307
rect 51771 106029 69493 106307
rect 69771 106029 87493 106307
rect 87771 106029 105493 106307
rect 105771 106029 123493 106307
rect 123771 106029 141493 106307
rect 141771 106029 159493 106307
rect 159771 106029 177493 106307
rect 177771 106029 195493 106307
rect 195771 106029 213493 106307
rect 213771 106029 231493 106307
rect 231771 106029 249493 106307
rect 249771 106029 267493 106307
rect 267771 106029 285493 106307
rect 285771 106029 296031 106307
rect 296309 106029 296325 106307
rect -4363 106013 296325 106029
rect -3403 104447 295365 104463
rect -3403 104169 -3387 104447
rect -3109 104169 13633 104447
rect 13911 104169 31633 104447
rect 31911 104169 49633 104447
rect 49911 104169 67633 104447
rect 67911 104169 85633 104447
rect 85911 104169 103633 104447
rect 103911 104169 121633 104447
rect 121911 104169 139633 104447
rect 139911 104169 157633 104447
rect 157911 104169 175633 104447
rect 175911 104169 193633 104447
rect 193911 104169 211633 104447
rect 211911 104169 229633 104447
rect 229911 104169 247633 104447
rect 247911 104169 265633 104447
rect 265911 104169 283633 104447
rect 283911 104169 295071 104447
rect 295349 104169 295365 104447
rect -3403 104153 295365 104169
rect -2443 102587 294405 102603
rect -2443 102309 -2427 102587
rect -2149 102309 11773 102587
rect 12051 102309 29773 102587
rect 30051 102309 47773 102587
rect 48051 102309 65773 102587
rect 66051 102309 83773 102587
rect 84051 102309 101773 102587
rect 102051 102309 119773 102587
rect 120051 102309 137773 102587
rect 138051 102309 155773 102587
rect 156051 102309 173773 102587
rect 174051 102309 191773 102587
rect 192051 102309 209773 102587
rect 210051 102309 227773 102587
rect 228051 102309 245773 102587
rect 246051 102309 263773 102587
rect 264051 102309 281773 102587
rect 282051 102309 294111 102587
rect 294389 102309 294405 102587
rect -2443 102293 294405 102309
rect -1483 100727 293445 100743
rect -1483 100449 -1467 100727
rect -1189 100449 9913 100727
rect 10191 100449 27913 100727
rect 28191 100449 45913 100727
rect 46191 100449 63913 100727
rect 64191 100449 81913 100727
rect 82191 100449 99913 100727
rect 100191 100449 117913 100727
rect 118191 100449 135913 100727
rect 136191 100449 153913 100727
rect 154191 100449 171913 100727
rect 172191 100449 189913 100727
rect 190191 100449 207913 100727
rect 208191 100449 225913 100727
rect 226191 100449 243913 100727
rect 244191 100449 261913 100727
rect 262191 100449 279913 100727
rect 280191 100449 293151 100727
rect 293429 100449 293445 100727
rect -1483 100433 293445 100449
rect -4363 97307 296325 97323
rect -4363 97029 -3867 97307
rect -3589 97029 6493 97307
rect 6771 97029 24493 97307
rect 24771 97029 42493 97307
rect 42771 97029 60493 97307
rect 60771 97029 78493 97307
rect 78771 97029 96493 97307
rect 96771 97029 114493 97307
rect 114771 97029 132493 97307
rect 132771 97029 150493 97307
rect 150771 97029 168493 97307
rect 168771 97029 186493 97307
rect 186771 97029 204493 97307
rect 204771 97029 222493 97307
rect 222771 97029 240493 97307
rect 240771 97029 258493 97307
rect 258771 97029 276493 97307
rect 276771 97029 295551 97307
rect 295829 97029 296325 97307
rect -4363 97013 296325 97029
rect -3403 95447 295365 95463
rect -3403 95169 -2907 95447
rect -2629 95169 4633 95447
rect 4911 95169 22633 95447
rect 22911 95169 40633 95447
rect 40911 95169 58633 95447
rect 58911 95169 76633 95447
rect 76911 95169 94633 95447
rect 94911 95169 112633 95447
rect 112911 95169 130633 95447
rect 130911 95169 148633 95447
rect 148911 95169 166633 95447
rect 166911 95169 184633 95447
rect 184911 95169 202633 95447
rect 202911 95169 220633 95447
rect 220911 95169 238633 95447
rect 238911 95169 256633 95447
rect 256911 95169 274633 95447
rect 274911 95169 294591 95447
rect 294869 95169 295365 95447
rect -3403 95153 295365 95169
rect -2443 93587 294405 93603
rect -2443 93309 -1947 93587
rect -1669 93309 2773 93587
rect 3051 93309 20773 93587
rect 21051 93309 38773 93587
rect 39051 93309 56773 93587
rect 57051 93309 74773 93587
rect 75051 93309 92773 93587
rect 93051 93309 110773 93587
rect 111051 93309 128773 93587
rect 129051 93309 146773 93587
rect 147051 93309 164773 93587
rect 165051 93309 182773 93587
rect 183051 93309 200773 93587
rect 201051 93309 218773 93587
rect 219051 93309 236773 93587
rect 237051 93309 254773 93587
rect 255051 93309 272773 93587
rect 273051 93309 290773 93587
rect 291051 93309 293631 93587
rect 293909 93309 294405 93587
rect -2443 93293 294405 93309
rect -1483 91727 293445 91743
rect -1483 91449 -987 91727
rect -709 91449 913 91727
rect 1191 91449 18913 91727
rect 19191 91449 36913 91727
rect 37191 91449 54913 91727
rect 55191 91449 72913 91727
rect 73191 91449 90913 91727
rect 91191 91449 108913 91727
rect 109191 91449 126913 91727
rect 127191 91449 144913 91727
rect 145191 91449 162913 91727
rect 163191 91449 180913 91727
rect 181191 91449 198913 91727
rect 199191 91449 216913 91727
rect 217191 91449 234913 91727
rect 235191 91449 252913 91727
rect 253191 91449 270913 91727
rect 271191 91449 288913 91727
rect 289191 91449 292671 91727
rect 292949 91449 293445 91727
rect -1483 91433 293445 91449
rect -4363 88307 296325 88323
rect -4363 88029 -4347 88307
rect -4069 88029 15493 88307
rect 15771 88029 33493 88307
rect 33771 88029 51493 88307
rect 51771 88029 69493 88307
rect 69771 88029 87493 88307
rect 87771 88029 105493 88307
rect 105771 88029 123493 88307
rect 123771 88029 141493 88307
rect 141771 88029 159493 88307
rect 159771 88029 177493 88307
rect 177771 88029 195493 88307
rect 195771 88029 213493 88307
rect 213771 88029 231493 88307
rect 231771 88029 249493 88307
rect 249771 88029 267493 88307
rect 267771 88029 285493 88307
rect 285771 88029 296031 88307
rect 296309 88029 296325 88307
rect -4363 88013 296325 88029
rect -3403 86447 295365 86463
rect -3403 86169 -3387 86447
rect -3109 86169 13633 86447
rect 13911 86169 31633 86447
rect 31911 86169 49633 86447
rect 49911 86169 67633 86447
rect 67911 86169 85633 86447
rect 85911 86169 103633 86447
rect 103911 86169 121633 86447
rect 121911 86169 139633 86447
rect 139911 86169 157633 86447
rect 157911 86169 175633 86447
rect 175911 86169 193633 86447
rect 193911 86169 211633 86447
rect 211911 86169 229633 86447
rect 229911 86169 247633 86447
rect 247911 86169 265633 86447
rect 265911 86169 283633 86447
rect 283911 86169 295071 86447
rect 295349 86169 295365 86447
rect -3403 86153 295365 86169
rect -2443 84587 294405 84603
rect -2443 84309 -2427 84587
rect -2149 84309 11773 84587
rect 12051 84309 29773 84587
rect 30051 84309 47773 84587
rect 48051 84309 65773 84587
rect 66051 84309 83773 84587
rect 84051 84309 101773 84587
rect 102051 84309 119773 84587
rect 120051 84309 137773 84587
rect 138051 84309 155773 84587
rect 156051 84309 173773 84587
rect 174051 84309 191773 84587
rect 192051 84309 209773 84587
rect 210051 84309 227773 84587
rect 228051 84309 245773 84587
rect 246051 84309 263773 84587
rect 264051 84309 281773 84587
rect 282051 84309 294111 84587
rect 294389 84309 294405 84587
rect -2443 84293 294405 84309
rect -1483 82727 293445 82743
rect -1483 82449 -1467 82727
rect -1189 82449 9913 82727
rect 10191 82449 27913 82727
rect 28191 82449 45913 82727
rect 46191 82449 63913 82727
rect 64191 82449 81913 82727
rect 82191 82449 99913 82727
rect 100191 82449 117913 82727
rect 118191 82449 135913 82727
rect 136191 82449 153913 82727
rect 154191 82449 171913 82727
rect 172191 82449 189913 82727
rect 190191 82449 207913 82727
rect 208191 82449 225913 82727
rect 226191 82449 243913 82727
rect 244191 82449 261913 82727
rect 262191 82449 279913 82727
rect 280191 82449 293151 82727
rect 293429 82449 293445 82727
rect -1483 82433 293445 82449
rect -4363 79307 296325 79323
rect -4363 79029 -3867 79307
rect -3589 79029 6493 79307
rect 6771 79029 24493 79307
rect 24771 79029 42493 79307
rect 42771 79029 60493 79307
rect 60771 79029 78493 79307
rect 78771 79029 96493 79307
rect 96771 79029 114493 79307
rect 114771 79029 132493 79307
rect 132771 79029 150493 79307
rect 150771 79029 168493 79307
rect 168771 79029 186493 79307
rect 186771 79029 204493 79307
rect 204771 79029 222493 79307
rect 222771 79029 240493 79307
rect 240771 79029 258493 79307
rect 258771 79029 276493 79307
rect 276771 79029 295551 79307
rect 295829 79029 296325 79307
rect -4363 79013 296325 79029
rect -3403 77447 295365 77463
rect -3403 77169 -2907 77447
rect -2629 77169 4633 77447
rect 4911 77169 22633 77447
rect 22911 77169 40633 77447
rect 40911 77169 58633 77447
rect 58911 77169 76633 77447
rect 76911 77169 94633 77447
rect 94911 77169 112633 77447
rect 112911 77169 130633 77447
rect 130911 77169 148633 77447
rect 148911 77169 166633 77447
rect 166911 77169 184633 77447
rect 184911 77169 202633 77447
rect 202911 77169 220633 77447
rect 220911 77169 238633 77447
rect 238911 77169 256633 77447
rect 256911 77169 274633 77447
rect 274911 77169 294591 77447
rect 294869 77169 295365 77447
rect -3403 77153 295365 77169
rect -2443 75587 294405 75603
rect -2443 75309 -1947 75587
rect -1669 75309 2773 75587
rect 3051 75309 20773 75587
rect 21051 75309 38773 75587
rect 39051 75309 56773 75587
rect 57051 75309 74773 75587
rect 75051 75309 92773 75587
rect 93051 75309 110773 75587
rect 111051 75309 128773 75587
rect 129051 75309 146773 75587
rect 147051 75309 164773 75587
rect 165051 75309 182773 75587
rect 183051 75309 200773 75587
rect 201051 75309 218773 75587
rect 219051 75309 236773 75587
rect 237051 75309 254773 75587
rect 255051 75309 272773 75587
rect 273051 75309 290773 75587
rect 291051 75309 293631 75587
rect 293909 75309 294405 75587
rect -2443 75293 294405 75309
rect -1483 73727 293445 73743
rect -1483 73449 -987 73727
rect -709 73449 913 73727
rect 1191 73449 18913 73727
rect 19191 73449 36913 73727
rect 37191 73449 54913 73727
rect 55191 73449 72913 73727
rect 73191 73449 90913 73727
rect 91191 73449 108913 73727
rect 109191 73449 126913 73727
rect 127191 73449 144913 73727
rect 145191 73449 162913 73727
rect 163191 73449 180913 73727
rect 181191 73449 198913 73727
rect 199191 73449 216913 73727
rect 217191 73449 234913 73727
rect 235191 73449 252913 73727
rect 253191 73449 270913 73727
rect 271191 73449 288913 73727
rect 289191 73449 292671 73727
rect 292949 73449 293445 73727
rect -1483 73433 293445 73449
rect -4363 70307 296325 70323
rect -4363 70029 -4347 70307
rect -4069 70029 15493 70307
rect 15771 70029 33493 70307
rect 33771 70029 51493 70307
rect 51771 70029 69493 70307
rect 69771 70029 87493 70307
rect 87771 70029 105493 70307
rect 105771 70029 123493 70307
rect 123771 70029 141493 70307
rect 141771 70029 159493 70307
rect 159771 70029 177493 70307
rect 177771 70029 195493 70307
rect 195771 70029 213493 70307
rect 213771 70029 231493 70307
rect 231771 70029 249493 70307
rect 249771 70029 267493 70307
rect 267771 70029 285493 70307
rect 285771 70029 296031 70307
rect 296309 70029 296325 70307
rect -4363 70013 296325 70029
rect -3403 68447 295365 68463
rect -3403 68169 -3387 68447
rect -3109 68169 13633 68447
rect 13911 68169 31633 68447
rect 31911 68169 49633 68447
rect 49911 68169 67633 68447
rect 67911 68169 85633 68447
rect 85911 68169 103633 68447
rect 103911 68169 121633 68447
rect 121911 68169 139633 68447
rect 139911 68169 157633 68447
rect 157911 68169 175633 68447
rect 175911 68169 193633 68447
rect 193911 68169 211633 68447
rect 211911 68169 229633 68447
rect 229911 68169 247633 68447
rect 247911 68169 265633 68447
rect 265911 68169 283633 68447
rect 283911 68169 295071 68447
rect 295349 68169 295365 68447
rect -3403 68153 295365 68169
rect -2443 66587 294405 66603
rect -2443 66309 -2427 66587
rect -2149 66309 11773 66587
rect 12051 66309 29773 66587
rect 30051 66309 47773 66587
rect 48051 66309 65773 66587
rect 66051 66309 83773 66587
rect 84051 66309 101773 66587
rect 102051 66309 119773 66587
rect 120051 66309 137773 66587
rect 138051 66309 155773 66587
rect 156051 66309 173773 66587
rect 174051 66309 191773 66587
rect 192051 66309 209773 66587
rect 210051 66309 227773 66587
rect 228051 66309 245773 66587
rect 246051 66309 263773 66587
rect 264051 66309 281773 66587
rect 282051 66309 294111 66587
rect 294389 66309 294405 66587
rect -2443 66293 294405 66309
rect -1483 64727 293445 64743
rect -1483 64449 -1467 64727
rect -1189 64449 9913 64727
rect 10191 64449 27913 64727
rect 28191 64449 45913 64727
rect 46191 64449 63913 64727
rect 64191 64449 81913 64727
rect 82191 64449 99913 64727
rect 100191 64449 117913 64727
rect 118191 64449 135913 64727
rect 136191 64449 153913 64727
rect 154191 64449 171913 64727
rect 172191 64449 189913 64727
rect 190191 64449 207913 64727
rect 208191 64449 225913 64727
rect 226191 64449 243913 64727
rect 244191 64449 261913 64727
rect 262191 64449 279913 64727
rect 280191 64449 293151 64727
rect 293429 64449 293445 64727
rect -1483 64433 293445 64449
rect -4363 61307 296325 61323
rect -4363 61029 -3867 61307
rect -3589 61029 6493 61307
rect 6771 61029 24493 61307
rect 24771 61029 42493 61307
rect 42771 61029 60493 61307
rect 60771 61029 78493 61307
rect 78771 61029 96493 61307
rect 96771 61029 114493 61307
rect 114771 61029 132493 61307
rect 132771 61029 150493 61307
rect 150771 61029 168493 61307
rect 168771 61029 186493 61307
rect 186771 61029 204493 61307
rect 204771 61029 222493 61307
rect 222771 61029 240493 61307
rect 240771 61029 258493 61307
rect 258771 61029 276493 61307
rect 276771 61029 295551 61307
rect 295829 61029 296325 61307
rect -4363 61013 296325 61029
rect -3403 59447 295365 59463
rect -3403 59169 -2907 59447
rect -2629 59169 4633 59447
rect 4911 59169 22633 59447
rect 22911 59169 40633 59447
rect 40911 59169 58633 59447
rect 58911 59169 76633 59447
rect 76911 59169 94633 59447
rect 94911 59169 112633 59447
rect 112911 59169 130633 59447
rect 130911 59169 148633 59447
rect 148911 59169 166633 59447
rect 166911 59169 184633 59447
rect 184911 59169 202633 59447
rect 202911 59169 220633 59447
rect 220911 59169 238633 59447
rect 238911 59169 256633 59447
rect 256911 59169 274633 59447
rect 274911 59169 294591 59447
rect 294869 59169 295365 59447
rect -3403 59153 295365 59169
rect -2443 57587 294405 57603
rect -2443 57309 -1947 57587
rect -1669 57309 2773 57587
rect 3051 57309 20773 57587
rect 21051 57309 38773 57587
rect 39051 57309 56773 57587
rect 57051 57309 74773 57587
rect 75051 57309 92773 57587
rect 93051 57309 110773 57587
rect 111051 57309 128773 57587
rect 129051 57309 146773 57587
rect 147051 57309 164773 57587
rect 165051 57309 182773 57587
rect 183051 57309 200773 57587
rect 201051 57309 218773 57587
rect 219051 57309 236773 57587
rect 237051 57309 254773 57587
rect 255051 57309 272773 57587
rect 273051 57309 290773 57587
rect 291051 57309 293631 57587
rect 293909 57309 294405 57587
rect -2443 57293 294405 57309
rect -1483 55727 293445 55743
rect -1483 55449 -987 55727
rect -709 55449 913 55727
rect 1191 55449 18913 55727
rect 19191 55449 36913 55727
rect 37191 55449 54913 55727
rect 55191 55449 72913 55727
rect 73191 55449 90913 55727
rect 91191 55449 108913 55727
rect 109191 55449 126913 55727
rect 127191 55449 144913 55727
rect 145191 55449 162913 55727
rect 163191 55449 180913 55727
rect 181191 55449 198913 55727
rect 199191 55449 216913 55727
rect 217191 55449 234913 55727
rect 235191 55449 252913 55727
rect 253191 55449 270913 55727
rect 271191 55449 288913 55727
rect 289191 55449 292671 55727
rect 292949 55449 293445 55727
rect -1483 55433 293445 55449
rect -4363 52307 296325 52323
rect -4363 52029 -4347 52307
rect -4069 52029 15493 52307
rect 15771 52029 33493 52307
rect 33771 52029 51493 52307
rect 51771 52029 69493 52307
rect 69771 52029 87493 52307
rect 87771 52029 105493 52307
rect 105771 52029 123493 52307
rect 123771 52029 141493 52307
rect 141771 52029 159493 52307
rect 159771 52029 177493 52307
rect 177771 52029 195493 52307
rect 195771 52029 213493 52307
rect 213771 52029 231493 52307
rect 231771 52029 249493 52307
rect 249771 52029 267493 52307
rect 267771 52029 285493 52307
rect 285771 52029 296031 52307
rect 296309 52029 296325 52307
rect -4363 52013 296325 52029
rect -3403 50447 295365 50463
rect -3403 50169 -3387 50447
rect -3109 50169 13633 50447
rect 13911 50169 31633 50447
rect 31911 50169 49633 50447
rect 49911 50169 67633 50447
rect 67911 50169 85633 50447
rect 85911 50169 103633 50447
rect 103911 50169 121633 50447
rect 121911 50169 139633 50447
rect 139911 50169 157633 50447
rect 157911 50169 175633 50447
rect 175911 50169 193633 50447
rect 193911 50169 211633 50447
rect 211911 50169 229633 50447
rect 229911 50169 247633 50447
rect 247911 50169 265633 50447
rect 265911 50169 283633 50447
rect 283911 50169 295071 50447
rect 295349 50169 295365 50447
rect -3403 50153 295365 50169
rect -2443 48587 294405 48603
rect -2443 48309 -2427 48587
rect -2149 48309 11773 48587
rect 12051 48309 29773 48587
rect 30051 48309 47773 48587
rect 48051 48309 65773 48587
rect 66051 48309 83773 48587
rect 84051 48309 101773 48587
rect 102051 48309 119773 48587
rect 120051 48309 137773 48587
rect 138051 48309 155773 48587
rect 156051 48309 173773 48587
rect 174051 48309 191773 48587
rect 192051 48309 209773 48587
rect 210051 48309 227773 48587
rect 228051 48309 245773 48587
rect 246051 48309 263773 48587
rect 264051 48309 281773 48587
rect 282051 48309 294111 48587
rect 294389 48309 294405 48587
rect -2443 48293 294405 48309
rect -1483 46727 293445 46743
rect -1483 46449 -1467 46727
rect -1189 46449 9913 46727
rect 10191 46449 27913 46727
rect 28191 46449 45913 46727
rect 46191 46449 63913 46727
rect 64191 46449 81913 46727
rect 82191 46449 99913 46727
rect 100191 46449 117913 46727
rect 118191 46449 135913 46727
rect 136191 46449 153913 46727
rect 154191 46449 171913 46727
rect 172191 46449 189913 46727
rect 190191 46449 207913 46727
rect 208191 46449 225913 46727
rect 226191 46449 243913 46727
rect 244191 46449 261913 46727
rect 262191 46449 279913 46727
rect 280191 46449 293151 46727
rect 293429 46449 293445 46727
rect -1483 46433 293445 46449
rect -4363 43307 296325 43323
rect -4363 43029 -3867 43307
rect -3589 43029 6493 43307
rect 6771 43029 24493 43307
rect 24771 43029 42493 43307
rect 42771 43029 60493 43307
rect 60771 43029 78493 43307
rect 78771 43029 96493 43307
rect 96771 43029 114493 43307
rect 114771 43029 132493 43307
rect 132771 43029 150493 43307
rect 150771 43029 168493 43307
rect 168771 43029 186493 43307
rect 186771 43029 204493 43307
rect 204771 43029 222493 43307
rect 222771 43029 240493 43307
rect 240771 43029 258493 43307
rect 258771 43029 276493 43307
rect 276771 43029 295551 43307
rect 295829 43029 296325 43307
rect -4363 43013 296325 43029
rect -3403 41447 295365 41463
rect -3403 41169 -2907 41447
rect -2629 41169 4633 41447
rect 4911 41169 22633 41447
rect 22911 41169 40633 41447
rect 40911 41169 58633 41447
rect 58911 41169 76633 41447
rect 76911 41169 94633 41447
rect 94911 41169 112633 41447
rect 112911 41169 130633 41447
rect 130911 41169 148633 41447
rect 148911 41169 166633 41447
rect 166911 41169 184633 41447
rect 184911 41169 202633 41447
rect 202911 41169 220633 41447
rect 220911 41169 238633 41447
rect 238911 41169 256633 41447
rect 256911 41169 274633 41447
rect 274911 41169 294591 41447
rect 294869 41169 295365 41447
rect -3403 41153 295365 41169
rect -2443 39587 294405 39603
rect -2443 39309 -1947 39587
rect -1669 39309 2773 39587
rect 3051 39309 20773 39587
rect 21051 39309 38773 39587
rect 39051 39309 56773 39587
rect 57051 39309 74773 39587
rect 75051 39309 92773 39587
rect 93051 39309 110773 39587
rect 111051 39309 128773 39587
rect 129051 39309 146773 39587
rect 147051 39309 164773 39587
rect 165051 39309 182773 39587
rect 183051 39309 200773 39587
rect 201051 39309 218773 39587
rect 219051 39309 236773 39587
rect 237051 39309 254773 39587
rect 255051 39309 272773 39587
rect 273051 39309 290773 39587
rect 291051 39309 293631 39587
rect 293909 39309 294405 39587
rect -2443 39293 294405 39309
rect -1483 37727 293445 37743
rect -1483 37449 -987 37727
rect -709 37449 913 37727
rect 1191 37449 18913 37727
rect 19191 37449 36913 37727
rect 37191 37449 54913 37727
rect 55191 37449 72913 37727
rect 73191 37449 90913 37727
rect 91191 37449 108913 37727
rect 109191 37449 126913 37727
rect 127191 37449 144913 37727
rect 145191 37449 162913 37727
rect 163191 37449 180913 37727
rect 181191 37449 198913 37727
rect 199191 37449 216913 37727
rect 217191 37449 234913 37727
rect 235191 37449 252913 37727
rect 253191 37449 270913 37727
rect 271191 37449 288913 37727
rect 289191 37449 292671 37727
rect 292949 37449 293445 37727
rect -1483 37433 293445 37449
rect -4363 34307 296325 34323
rect -4363 34029 -4347 34307
rect -4069 34029 15493 34307
rect 15771 34029 33493 34307
rect 33771 34029 51493 34307
rect 51771 34029 69493 34307
rect 69771 34029 87493 34307
rect 87771 34029 105493 34307
rect 105771 34029 123493 34307
rect 123771 34029 141493 34307
rect 141771 34029 159493 34307
rect 159771 34029 177493 34307
rect 177771 34029 195493 34307
rect 195771 34029 213493 34307
rect 213771 34029 231493 34307
rect 231771 34029 249493 34307
rect 249771 34029 267493 34307
rect 267771 34029 285493 34307
rect 285771 34029 296031 34307
rect 296309 34029 296325 34307
rect -4363 34013 296325 34029
rect -3403 32447 295365 32463
rect -3403 32169 -3387 32447
rect -3109 32169 13633 32447
rect 13911 32169 31633 32447
rect 31911 32169 49633 32447
rect 49911 32169 67633 32447
rect 67911 32169 85633 32447
rect 85911 32169 103633 32447
rect 103911 32169 121633 32447
rect 121911 32169 139633 32447
rect 139911 32169 157633 32447
rect 157911 32169 175633 32447
rect 175911 32169 193633 32447
rect 193911 32169 211633 32447
rect 211911 32169 229633 32447
rect 229911 32169 247633 32447
rect 247911 32169 265633 32447
rect 265911 32169 283633 32447
rect 283911 32169 295071 32447
rect 295349 32169 295365 32447
rect -3403 32153 295365 32169
rect -2443 30587 294405 30603
rect -2443 30309 -2427 30587
rect -2149 30309 11773 30587
rect 12051 30309 29773 30587
rect 30051 30309 47773 30587
rect 48051 30309 65773 30587
rect 66051 30309 83773 30587
rect 84051 30309 101773 30587
rect 102051 30309 119773 30587
rect 120051 30309 137773 30587
rect 138051 30309 155773 30587
rect 156051 30309 173773 30587
rect 174051 30309 191773 30587
rect 192051 30309 209773 30587
rect 210051 30309 227773 30587
rect 228051 30309 245773 30587
rect 246051 30309 263773 30587
rect 264051 30309 281773 30587
rect 282051 30309 294111 30587
rect 294389 30309 294405 30587
rect -2443 30293 294405 30309
rect -1483 28727 293445 28743
rect -1483 28449 -1467 28727
rect -1189 28449 9913 28727
rect 10191 28449 27913 28727
rect 28191 28449 45913 28727
rect 46191 28449 63913 28727
rect 64191 28449 81913 28727
rect 82191 28449 99913 28727
rect 100191 28449 117913 28727
rect 118191 28449 135913 28727
rect 136191 28449 153913 28727
rect 154191 28449 171913 28727
rect 172191 28449 189913 28727
rect 190191 28449 207913 28727
rect 208191 28449 225913 28727
rect 226191 28449 243913 28727
rect 244191 28449 261913 28727
rect 262191 28449 279913 28727
rect 280191 28449 293151 28727
rect 293429 28449 293445 28727
rect -1483 28433 293445 28449
rect -4363 25307 296325 25323
rect -4363 25029 -3867 25307
rect -3589 25029 6493 25307
rect 6771 25029 24493 25307
rect 24771 25029 42493 25307
rect 42771 25029 60493 25307
rect 60771 25029 78493 25307
rect 78771 25029 96493 25307
rect 96771 25029 114493 25307
rect 114771 25029 132493 25307
rect 132771 25029 150493 25307
rect 150771 25029 168493 25307
rect 168771 25029 186493 25307
rect 186771 25029 204493 25307
rect 204771 25029 222493 25307
rect 222771 25029 240493 25307
rect 240771 25029 258493 25307
rect 258771 25029 276493 25307
rect 276771 25029 295551 25307
rect 295829 25029 296325 25307
rect -4363 25013 296325 25029
rect -3403 23447 295365 23463
rect -3403 23169 -2907 23447
rect -2629 23169 4633 23447
rect 4911 23169 22633 23447
rect 22911 23169 40633 23447
rect 40911 23169 58633 23447
rect 58911 23169 76633 23447
rect 76911 23169 94633 23447
rect 94911 23169 112633 23447
rect 112911 23169 130633 23447
rect 130911 23169 148633 23447
rect 148911 23169 166633 23447
rect 166911 23169 184633 23447
rect 184911 23169 202633 23447
rect 202911 23169 220633 23447
rect 220911 23169 238633 23447
rect 238911 23169 256633 23447
rect 256911 23169 274633 23447
rect 274911 23169 294591 23447
rect 294869 23169 295365 23447
rect -3403 23153 295365 23169
rect -2443 21587 294405 21603
rect -2443 21309 -1947 21587
rect -1669 21309 2773 21587
rect 3051 21309 20773 21587
rect 21051 21309 38773 21587
rect 39051 21309 56773 21587
rect 57051 21309 74773 21587
rect 75051 21309 92773 21587
rect 93051 21309 110773 21587
rect 111051 21309 128773 21587
rect 129051 21309 146773 21587
rect 147051 21309 164773 21587
rect 165051 21309 182773 21587
rect 183051 21309 200773 21587
rect 201051 21309 218773 21587
rect 219051 21309 236773 21587
rect 237051 21309 254773 21587
rect 255051 21309 272773 21587
rect 273051 21309 290773 21587
rect 291051 21309 293631 21587
rect 293909 21309 294405 21587
rect -2443 21293 294405 21309
rect -1483 19727 293445 19743
rect -1483 19449 -987 19727
rect -709 19449 913 19727
rect 1191 19449 18913 19727
rect 19191 19449 36913 19727
rect 37191 19449 54913 19727
rect 55191 19449 72913 19727
rect 73191 19449 90913 19727
rect 91191 19449 108913 19727
rect 109191 19449 126913 19727
rect 127191 19449 144913 19727
rect 145191 19449 162913 19727
rect 163191 19449 180913 19727
rect 181191 19449 198913 19727
rect 199191 19449 216913 19727
rect 217191 19449 234913 19727
rect 235191 19449 252913 19727
rect 253191 19449 270913 19727
rect 271191 19449 288913 19727
rect 289191 19449 292671 19727
rect 292949 19449 293445 19727
rect -1483 19433 293445 19449
rect -4363 16307 296325 16323
rect -4363 16029 -4347 16307
rect -4069 16029 15493 16307
rect 15771 16029 33493 16307
rect 33771 16029 51493 16307
rect 51771 16029 69493 16307
rect 69771 16029 87493 16307
rect 87771 16029 105493 16307
rect 105771 16029 123493 16307
rect 123771 16029 141493 16307
rect 141771 16029 159493 16307
rect 159771 16029 177493 16307
rect 177771 16029 195493 16307
rect 195771 16029 213493 16307
rect 213771 16029 231493 16307
rect 231771 16029 249493 16307
rect 249771 16029 267493 16307
rect 267771 16029 285493 16307
rect 285771 16029 296031 16307
rect 296309 16029 296325 16307
rect -4363 16013 296325 16029
rect -3403 14447 295365 14463
rect -3403 14169 -3387 14447
rect -3109 14169 13633 14447
rect 13911 14169 31633 14447
rect 31911 14169 49633 14447
rect 49911 14169 67633 14447
rect 67911 14169 85633 14447
rect 85911 14169 103633 14447
rect 103911 14169 121633 14447
rect 121911 14169 139633 14447
rect 139911 14169 157633 14447
rect 157911 14169 175633 14447
rect 175911 14169 193633 14447
rect 193911 14169 211633 14447
rect 211911 14169 229633 14447
rect 229911 14169 247633 14447
rect 247911 14169 265633 14447
rect 265911 14169 283633 14447
rect 283911 14169 295071 14447
rect 295349 14169 295365 14447
rect -3403 14153 295365 14169
rect -2443 12587 294405 12603
rect -2443 12309 -2427 12587
rect -2149 12309 11773 12587
rect 12051 12309 29773 12587
rect 30051 12309 47773 12587
rect 48051 12309 65773 12587
rect 66051 12309 83773 12587
rect 84051 12309 101773 12587
rect 102051 12309 119773 12587
rect 120051 12309 137773 12587
rect 138051 12309 155773 12587
rect 156051 12309 173773 12587
rect 174051 12309 191773 12587
rect 192051 12309 209773 12587
rect 210051 12309 227773 12587
rect 228051 12309 245773 12587
rect 246051 12309 263773 12587
rect 264051 12309 281773 12587
rect 282051 12309 294111 12587
rect 294389 12309 294405 12587
rect -2443 12293 294405 12309
rect -1483 10727 293445 10743
rect -1483 10449 -1467 10727
rect -1189 10449 9913 10727
rect 10191 10449 27913 10727
rect 28191 10449 45913 10727
rect 46191 10449 63913 10727
rect 64191 10449 81913 10727
rect 82191 10449 99913 10727
rect 100191 10449 117913 10727
rect 118191 10449 135913 10727
rect 136191 10449 153913 10727
rect 154191 10449 171913 10727
rect 172191 10449 189913 10727
rect 190191 10449 207913 10727
rect 208191 10449 225913 10727
rect 226191 10449 243913 10727
rect 244191 10449 261913 10727
rect 262191 10449 279913 10727
rect 280191 10449 293151 10727
rect 293429 10449 293445 10727
rect -1483 10433 293445 10449
rect -4363 7307 296325 7323
rect -4363 7029 -3867 7307
rect -3589 7029 6493 7307
rect 6771 7029 24493 7307
rect 24771 7029 42493 7307
rect 42771 7029 60493 7307
rect 60771 7029 78493 7307
rect 78771 7029 96493 7307
rect 96771 7029 114493 7307
rect 114771 7029 132493 7307
rect 132771 7029 150493 7307
rect 150771 7029 168493 7307
rect 168771 7029 186493 7307
rect 186771 7029 204493 7307
rect 204771 7029 222493 7307
rect 222771 7029 240493 7307
rect 240771 7029 258493 7307
rect 258771 7029 276493 7307
rect 276771 7029 295551 7307
rect 295829 7029 296325 7307
rect -4363 7013 296325 7029
rect -3403 5447 295365 5463
rect -3403 5169 -2907 5447
rect -2629 5169 4633 5447
rect 4911 5169 22633 5447
rect 22911 5169 40633 5447
rect 40911 5169 58633 5447
rect 58911 5169 76633 5447
rect 76911 5169 94633 5447
rect 94911 5169 112633 5447
rect 112911 5169 130633 5447
rect 130911 5169 148633 5447
rect 148911 5169 166633 5447
rect 166911 5169 184633 5447
rect 184911 5169 202633 5447
rect 202911 5169 220633 5447
rect 220911 5169 238633 5447
rect 238911 5169 256633 5447
rect 256911 5169 274633 5447
rect 274911 5169 294591 5447
rect 294869 5169 295365 5447
rect -3403 5153 295365 5169
rect -2443 3587 294405 3603
rect -2443 3309 -1947 3587
rect -1669 3309 2773 3587
rect 3051 3309 20773 3587
rect 21051 3309 38773 3587
rect 39051 3309 56773 3587
rect 57051 3309 74773 3587
rect 75051 3309 92773 3587
rect 93051 3309 110773 3587
rect 111051 3309 128773 3587
rect 129051 3309 146773 3587
rect 147051 3309 164773 3587
rect 165051 3309 182773 3587
rect 183051 3309 200773 3587
rect 201051 3309 218773 3587
rect 219051 3309 236773 3587
rect 237051 3309 254773 3587
rect 255051 3309 272773 3587
rect 273051 3309 290773 3587
rect 291051 3309 293631 3587
rect 293909 3309 294405 3587
rect -2443 3293 294405 3309
rect -1483 1727 293445 1743
rect -1483 1449 -987 1727
rect -709 1449 913 1727
rect 1191 1449 18913 1727
rect 19191 1449 36913 1727
rect 37191 1449 54913 1727
rect 55191 1449 72913 1727
rect 73191 1449 90913 1727
rect 91191 1449 108913 1727
rect 109191 1449 126913 1727
rect 127191 1449 144913 1727
rect 145191 1449 162913 1727
rect 163191 1449 180913 1727
rect 181191 1449 198913 1727
rect 199191 1449 216913 1727
rect 217191 1449 234913 1727
rect 235191 1449 252913 1727
rect 253191 1449 270913 1727
rect 271191 1449 288913 1727
rect 289191 1449 292671 1727
rect 292949 1449 293445 1727
rect -1483 1433 293445 1449
rect -1003 -173 292965 -157
rect -1003 -451 -987 -173
rect -709 -451 913 -173
rect 1191 -451 18913 -173
rect 19191 -451 36913 -173
rect 37191 -451 54913 -173
rect 55191 -451 72913 -173
rect 73191 -451 90913 -173
rect 91191 -451 108913 -173
rect 109191 -451 126913 -173
rect 127191 -451 144913 -173
rect 145191 -451 162913 -173
rect 163191 -451 180913 -173
rect 181191 -451 198913 -173
rect 199191 -451 216913 -173
rect 217191 -451 234913 -173
rect 235191 -451 252913 -173
rect 253191 -451 270913 -173
rect 271191 -451 288913 -173
rect 289191 -451 292671 -173
rect 292949 -451 292965 -173
rect -1003 -467 292965 -451
rect -1483 -653 293445 -637
rect -1483 -931 -1467 -653
rect -1189 -931 9913 -653
rect 10191 -931 27913 -653
rect 28191 -931 45913 -653
rect 46191 -931 63913 -653
rect 64191 -931 81913 -653
rect 82191 -931 99913 -653
rect 100191 -931 117913 -653
rect 118191 -931 135913 -653
rect 136191 -931 153913 -653
rect 154191 -931 171913 -653
rect 172191 -931 189913 -653
rect 190191 -931 207913 -653
rect 208191 -931 225913 -653
rect 226191 -931 243913 -653
rect 244191 -931 261913 -653
rect 262191 -931 279913 -653
rect 280191 -931 293151 -653
rect 293429 -931 293445 -653
rect -1483 -947 293445 -931
rect -1963 -1133 293925 -1117
rect -1963 -1411 -1947 -1133
rect -1669 -1411 2773 -1133
rect 3051 -1411 20773 -1133
rect 21051 -1411 38773 -1133
rect 39051 -1411 56773 -1133
rect 57051 -1411 74773 -1133
rect 75051 -1411 92773 -1133
rect 93051 -1411 110773 -1133
rect 111051 -1411 128773 -1133
rect 129051 -1411 146773 -1133
rect 147051 -1411 164773 -1133
rect 165051 -1411 182773 -1133
rect 183051 -1411 200773 -1133
rect 201051 -1411 218773 -1133
rect 219051 -1411 236773 -1133
rect 237051 -1411 254773 -1133
rect 255051 -1411 272773 -1133
rect 273051 -1411 290773 -1133
rect 291051 -1411 293631 -1133
rect 293909 -1411 293925 -1133
rect -1963 -1427 293925 -1411
rect -2443 -1613 294405 -1597
rect -2443 -1891 -2427 -1613
rect -2149 -1891 11773 -1613
rect 12051 -1891 29773 -1613
rect 30051 -1891 47773 -1613
rect 48051 -1891 65773 -1613
rect 66051 -1891 83773 -1613
rect 84051 -1891 101773 -1613
rect 102051 -1891 119773 -1613
rect 120051 -1891 137773 -1613
rect 138051 -1891 155773 -1613
rect 156051 -1891 173773 -1613
rect 174051 -1891 191773 -1613
rect 192051 -1891 209773 -1613
rect 210051 -1891 227773 -1613
rect 228051 -1891 245773 -1613
rect 246051 -1891 263773 -1613
rect 264051 -1891 281773 -1613
rect 282051 -1891 294111 -1613
rect 294389 -1891 294405 -1613
rect -2443 -1907 294405 -1891
rect -2923 -2093 294885 -2077
rect -2923 -2371 -2907 -2093
rect -2629 -2371 4633 -2093
rect 4911 -2371 22633 -2093
rect 22911 -2371 40633 -2093
rect 40911 -2371 58633 -2093
rect 58911 -2371 76633 -2093
rect 76911 -2371 94633 -2093
rect 94911 -2371 112633 -2093
rect 112911 -2371 130633 -2093
rect 130911 -2371 148633 -2093
rect 148911 -2371 166633 -2093
rect 166911 -2371 184633 -2093
rect 184911 -2371 202633 -2093
rect 202911 -2371 220633 -2093
rect 220911 -2371 238633 -2093
rect 238911 -2371 256633 -2093
rect 256911 -2371 274633 -2093
rect 274911 -2371 294591 -2093
rect 294869 -2371 294885 -2093
rect -2923 -2387 294885 -2371
rect -3403 -2573 295365 -2557
rect -3403 -2851 -3387 -2573
rect -3109 -2851 13633 -2573
rect 13911 -2851 31633 -2573
rect 31911 -2851 49633 -2573
rect 49911 -2851 67633 -2573
rect 67911 -2851 85633 -2573
rect 85911 -2851 103633 -2573
rect 103911 -2851 121633 -2573
rect 121911 -2851 139633 -2573
rect 139911 -2851 157633 -2573
rect 157911 -2851 175633 -2573
rect 175911 -2851 193633 -2573
rect 193911 -2851 211633 -2573
rect 211911 -2851 229633 -2573
rect 229911 -2851 247633 -2573
rect 247911 -2851 265633 -2573
rect 265911 -2851 283633 -2573
rect 283911 -2851 295071 -2573
rect 295349 -2851 295365 -2573
rect -3403 -2867 295365 -2851
rect -3883 -3053 295845 -3037
rect -3883 -3331 -3867 -3053
rect -3589 -3331 6493 -3053
rect 6771 -3331 24493 -3053
rect 24771 -3331 42493 -3053
rect 42771 -3331 60493 -3053
rect 60771 -3331 78493 -3053
rect 78771 -3331 96493 -3053
rect 96771 -3331 114493 -3053
rect 114771 -3331 132493 -3053
rect 132771 -3331 150493 -3053
rect 150771 -3331 168493 -3053
rect 168771 -3331 186493 -3053
rect 186771 -3331 204493 -3053
rect 204771 -3331 222493 -3053
rect 222771 -3331 240493 -3053
rect 240771 -3331 258493 -3053
rect 258771 -3331 276493 -3053
rect 276771 -3331 295551 -3053
rect 295829 -3331 295845 -3053
rect -3883 -3347 295845 -3331
rect -4363 -3533 296325 -3517
rect -4363 -3811 -4347 -3533
rect -4069 -3811 15493 -3533
rect 15771 -3811 33493 -3533
rect 33771 -3811 51493 -3533
rect 51771 -3811 69493 -3533
rect 69771 -3811 87493 -3533
rect 87771 -3811 105493 -3533
rect 105771 -3811 123493 -3533
rect 123771 -3811 141493 -3533
rect 141771 -3811 159493 -3533
rect 159771 -3811 177493 -3533
rect 177771 -3811 195493 -3533
rect 195771 -3811 213493 -3533
rect 213771 -3811 231493 -3533
rect 231771 -3811 249493 -3533
rect 249771 -3811 267493 -3533
rect 267771 -3811 285493 -3533
rect 285771 -3811 296031 -3533
rect 296309 -3811 296325 -3533
rect -4363 -3827 296325 -3811
<< labels >>
rlabel metal3 s 291760 142638 292480 142758 4 analog_io[0]
port 1 nsew
rlabel metal2 s 223049 351760 223105 352480 4 analog_io[10]
port 2 nsew
rlabel metal2 s 190573 351760 190629 352480 4 analog_io[11]
port 3 nsew
rlabel metal2 s 158143 351760 158199 352480 4 analog_io[12]
port 4 nsew
rlabel metal2 s 125713 351760 125769 352480 4 analog_io[13]
port 5 nsew
rlabel metal2 s 93237 351760 93293 352480 4 analog_io[14]
port 6 nsew
rlabel metal2 s 60807 351760 60863 352480 4 analog_io[15]
port 7 nsew
rlabel metal2 s 28377 351760 28433 352480 4 analog_io[16]
port 8 nsew
rlabel metal3 s -480 348610 240 348730 4 analog_io[17]
port 9 nsew
rlabel metal3 s -480 322498 240 322618 4 analog_io[18]
port 10 nsew
rlabel metal3 s -480 296454 240 296574 4 analog_io[19]
port 11 nsew
rlabel metal3 s 291760 169226 292480 169346 4 analog_io[1]
port 12 nsew
rlabel metal3 s -480 270342 240 270462 4 analog_io[20]
port 13 nsew
rlabel metal3 s -480 244298 240 244418 4 analog_io[21]
port 14 nsew
rlabel metal3 s -480 218254 240 218374 4 analog_io[22]
port 15 nsew
rlabel metal3 s -480 192142 240 192262 4 analog_io[23]
port 16 nsew
rlabel metal3 s -480 166098 240 166218 4 analog_io[24]
port 17 nsew
rlabel metal3 s -480 139986 240 140106 4 analog_io[25]
port 18 nsew
rlabel metal3 s -480 113942 240 114062 4 analog_io[26]
port 19 nsew
rlabel metal3 s -480 87898 240 88018 4 analog_io[27]
port 20 nsew
rlabel metal3 s -480 61786 240 61906 4 analog_io[28]
port 21 nsew
rlabel metal3 s 291760 195814 292480 195934 4 analog_io[2]
port 22 nsew
rlabel metal3 s 291760 222334 292480 222454 4 analog_io[3]
port 23 nsew
rlabel metal3 s 291760 248922 292480 249042 4 analog_io[4]
port 24 nsew
rlabel metal3 s 291760 275510 292480 275630 4 analog_io[5]
port 25 nsew
rlabel metal3 s 291760 302030 292480 302150 4 analog_io[6]
port 26 nsew
rlabel metal3 s 291760 328618 292480 328738 4 analog_io[7]
port 27 nsew
rlabel metal2 s 287909 351760 287965 352480 4 analog_io[8]
port 28 nsew
rlabel metal2 s 255479 351760 255535 352480 4 analog_io[9]
port 29 nsew
rlabel metal3 s 291760 3238 292480 3358 4 io_in[0]
port 30 nsew
rlabel metal3 s 291760 9834 292480 9954 4 io_out[0]
port 31 nsew
rlabel metal3 s 291760 228998 292480 229118 4 io_in[10]
port 32 nsew
rlabel metal3 s 291760 235662 292480 235782 4 io_out[10]
port 33 nsew
rlabel metal3 s 291760 255586 292480 255706 4 io_in[11]
port 34 nsew
rlabel metal3 s 291760 262182 292480 262302 4 io_out[11]
port 35 nsew
rlabel metal3 s 291760 282106 292480 282226 4 io_in[12]
port 36 nsew
rlabel metal3 s 291760 288770 292480 288890 4 io_out[12]
port 37 nsew
rlabel metal3 s 291760 308694 292480 308814 4 io_in[13]
port 38 nsew
rlabel metal3 s 291760 315358 292480 315478 4 io_out[13]
port 39 nsew
rlabel metal3 s 291760 335282 292480 335402 4 io_in[14]
port 40 nsew
rlabel metal3 s 291760 341878 292480 341998 4 io_out[14]
port 41 nsew
rlabel metal2 s 279813 351760 279869 352480 4 io_in[15]
port 42 nsew
rlabel metal2 s 271717 351760 271773 352480 4 io_out[15]
port 43 nsew
rlabel metal2 s 247383 351760 247439 352480 4 io_in[16]
port 44 nsew
rlabel metal2 s 239241 351760 239297 352480 4 io_out[16]
port 45 nsew
rlabel metal2 s 214907 351760 214963 352480 4 io_in[17]
port 46 nsew
rlabel metal2 s 206811 351760 206867 352480 4 io_out[17]
port 47 nsew
rlabel metal2 s 182477 351760 182533 352480 4 io_in[18]
port 48 nsew
rlabel metal2 s 174381 351760 174437 352480 4 io_out[18]
port 49 nsew
rlabel metal2 s 150047 351760 150103 352480 4 io_in[19]
port 50 nsew
rlabel metal2 s 141905 351760 141961 352480 4 io_out[19]
port 51 nsew
rlabel metal3 s 291760 23094 292480 23214 4 io_in[1]
port 52 nsew
rlabel metal3 s 291760 29758 292480 29878 4 io_out[1]
port 53 nsew
rlabel metal2 s 117571 351760 117627 352480 4 io_in[20]
port 54 nsew
rlabel metal2 s 109475 351760 109531 352480 4 io_out[20]
port 55 nsew
rlabel metal2 s 85141 351760 85197 352480 4 io_in[21]
port 56 nsew
rlabel metal2 s 77045 351760 77101 352480 4 io_out[21]
port 57 nsew
rlabel metal2 s 52711 351760 52767 352480 4 io_in[22]
port 58 nsew
rlabel metal2 s 44569 351760 44625 352480 4 io_out[22]
port 59 nsew
rlabel metal2 s 20235 351760 20291 352480 4 io_in[23]
port 60 nsew
rlabel metal2 s 12139 351760 12195 352480 4 io_out[23]
port 61 nsew
rlabel metal3 s -480 342082 240 342202 4 io_in[24]
port 62 nsew
rlabel metal3 s -480 335554 240 335674 4 io_out[24]
port 63 nsew
rlabel metal3 s -480 315970 240 316090 4 io_in[25]
port 64 nsew
rlabel metal3 s -480 309510 240 309630 4 io_out[25]
port 65 nsew
rlabel metal3 s -480 289926 240 290046 4 io_in[26]
port 66 nsew
rlabel metal3 s -480 283398 240 283518 4 io_out[26]
port 67 nsew
rlabel metal3 s -480 263882 240 264002 4 io_in[27]
port 68 nsew
rlabel metal3 s -480 257354 240 257474 4 io_out[27]
port 69 nsew
rlabel metal3 s -480 237770 240 237890 4 io_in[28]
port 70 nsew
rlabel metal3 s -480 231242 240 231362 4 io_out[28]
port 71 nsew
rlabel metal3 s -480 211726 240 211846 4 io_in[29]
port 72 nsew
rlabel metal3 s -480 205198 240 205318 4 io_out[29]
port 73 nsew
rlabel metal3 s 291760 43018 292480 43138 4 io_in[2]
port 74 nsew
rlabel metal3 s 291760 49682 292480 49802 4 io_out[2]
port 75 nsew
rlabel metal3 s -480 185614 240 185734 4 io_in[30]
port 76 nsew
rlabel metal3 s -480 179154 240 179274 4 io_out[30]
port 77 nsew
rlabel metal3 s -480 159570 240 159690 4 io_in[31]
port 78 nsew
rlabel metal3 s -480 153042 240 153162 4 io_out[31]
port 79 nsew
rlabel metal3 s -480 133526 240 133646 4 io_in[32]
port 80 nsew
rlabel metal3 s -480 126998 240 127118 4 io_out[32]
port 81 nsew
rlabel metal3 s -480 107414 240 107534 4 io_in[33]
port 82 nsew
rlabel metal3 s -480 100886 240 101006 4 io_out[33]
port 83 nsew
rlabel metal3 s -480 81370 240 81490 4 io_in[34]
port 84 nsew
rlabel metal3 s -480 74842 240 74962 4 io_out[34]
port 85 nsew
rlabel metal3 s -480 55258 240 55378 4 io_in[35]
port 86 nsew
rlabel metal3 s -480 48730 240 48850 4 io_out[35]
port 87 nsew
rlabel metal3 s -480 35742 240 35862 4 io_in[36]
port 88 nsew
rlabel metal3 s -480 29214 240 29334 4 io_out[36]
port 89 nsew
rlabel metal3 s -480 16158 240 16278 4 io_in[37]
port 90 nsew
rlabel metal3 s -480 9630 240 9750 4 io_out[37]
port 91 nsew
rlabel metal3 s 291760 62942 292480 63062 4 io_in[3]
port 92 nsew
rlabel metal3 s 291760 69606 292480 69726 4 io_out[3]
port 93 nsew
rlabel metal3 s 291760 82866 292480 82986 4 io_in[4]
port 94 nsew
rlabel metal3 s 291760 89530 292480 89650 4 io_out[4]
port 95 nsew
rlabel metal3 s 291760 102790 292480 102910 4 io_in[5]
port 96 nsew
rlabel metal3 s 291760 109454 292480 109574 4 io_out[5]
port 97 nsew
rlabel metal3 s 291760 122714 292480 122834 4 io_in[6]
port 98 nsew
rlabel metal3 s 291760 129378 292480 129498 4 io_out[6]
port 99 nsew
rlabel metal3 s 291760 149302 292480 149422 4 io_in[7]
port 100 nsew
rlabel metal3 s 291760 155966 292480 156086 4 io_out[7]
port 101 nsew
rlabel metal3 s 291760 175890 292480 176010 4 io_in[8]
port 102 nsew
rlabel metal3 s 291760 182486 292480 182606 4 io_out[8]
port 103 nsew
rlabel metal3 s 291760 202410 292480 202530 4 io_in[9]
port 104 nsew
rlabel metal3 s 291760 209074 292480 209194 4 io_out[9]
port 105 nsew
rlabel metal3 s 291760 16498 292480 16618 4 io_oeb[0]
port 106 nsew
rlabel metal3 s 291760 242258 292480 242378 4 io_oeb[10]
port 107 nsew
rlabel metal3 s 291760 268846 292480 268966 4 io_oeb[11]
port 108 nsew
rlabel metal3 s 291760 295434 292480 295554 4 io_oeb[12]
port 109 nsew
rlabel metal3 s 291760 321954 292480 322074 4 io_oeb[13]
port 110 nsew
rlabel metal3 s 291760 348542 292480 348662 4 io_oeb[14]
port 111 nsew
rlabel metal2 s 263575 351760 263631 352480 4 io_oeb[15]
port 112 nsew
rlabel metal2 s 231145 351760 231201 352480 4 io_oeb[16]
port 113 nsew
rlabel metal2 s 198715 351760 198771 352480 4 io_oeb[17]
port 114 nsew
rlabel metal2 s 166239 351760 166295 352480 4 io_oeb[18]
port 115 nsew
rlabel metal2 s 133809 351760 133865 352480 4 io_oeb[19]
port 116 nsew
rlabel metal3 s 291760 36422 292480 36542 4 io_oeb[1]
port 117 nsew
rlabel metal2 s 101379 351760 101435 352480 4 io_oeb[20]
port 118 nsew
rlabel metal2 s 68903 351760 68959 352480 4 io_oeb[21]
port 119 nsew
rlabel metal2 s 36473 351760 36529 352480 4 io_oeb[22]
port 120 nsew
rlabel metal2 s 4043 351760 4099 352480 4 io_oeb[23]
port 121 nsew
rlabel metal3 s -480 329026 240 329146 4 io_oeb[24]
port 122 nsew
rlabel metal3 s -480 302982 240 303102 4 io_oeb[25]
port 123 nsew
rlabel metal3 s -480 276870 240 276990 4 io_oeb[26]
port 124 nsew
rlabel metal3 s -480 250826 240 250946 4 io_oeb[27]
port 125 nsew
rlabel metal3 s -480 224714 240 224834 4 io_oeb[28]
port 126 nsew
rlabel metal3 s -480 198670 240 198790 4 io_oeb[29]
port 127 nsew
rlabel metal3 s 291760 56346 292480 56466 4 io_oeb[2]
port 128 nsew
rlabel metal3 s -480 172626 240 172746 4 io_oeb[30]
port 129 nsew
rlabel metal3 s -480 146514 240 146634 4 io_oeb[31]
port 130 nsew
rlabel metal3 s -480 120470 240 120590 4 io_oeb[32]
port 131 nsew
rlabel metal3 s -480 94358 240 94478 4 io_oeb[33]
port 132 nsew
rlabel metal3 s -480 68314 240 68434 4 io_oeb[34]
port 133 nsew
rlabel metal3 s -480 42270 240 42390 4 io_oeb[35]
port 134 nsew
rlabel metal3 s -480 22686 240 22806 4 io_oeb[36]
port 135 nsew
rlabel metal3 s -480 3170 240 3290 4 io_oeb[37]
port 136 nsew
rlabel metal3 s 291760 76270 292480 76390 4 io_oeb[3]
port 137 nsew
rlabel metal3 s 291760 96194 292480 96314 4 io_oeb[4]
port 138 nsew
rlabel metal3 s 291760 116118 292480 116238 4 io_oeb[5]
port 139 nsew
rlabel metal3 s 291760 136042 292480 136162 4 io_oeb[6]
port 140 nsew
rlabel metal3 s 291760 162562 292480 162682 4 io_oeb[7]
port 141 nsew
rlabel metal3 s 291760 189150 292480 189270 4 io_oeb[8]
port 142 nsew
rlabel metal3 s 291760 215738 292480 215858 4 io_oeb[9]
port 143 nsew
rlabel metal2 s 62923 -480 62979 240 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 240253 -480 240309 240 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 242001 -480 242057 240 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 243795 -480 243851 240 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 245543 -480 245599 240 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 247337 -480 247393 240 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 249085 -480 249141 240 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 250879 -480 250935 240 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 252673 -480 252729 240 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 254421 -480 254477 240 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 256215 -480 256271 240 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 80633 -480 80689 240 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 257963 -480 258019 240 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 259757 -480 259813 240 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 261505 -480 261561 240 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 263299 -480 263355 240 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 265047 -480 265103 240 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 266841 -480 266897 240 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 268589 -480 268645 240 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 270383 -480 270439 240 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 272177 -480 272233 240 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 273925 -480 273981 240 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 82427 -480 82483 240 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 275719 -480 275775 240 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 277467 -480 277523 240 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 279261 -480 279317 240 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 281009 -480 281065 240 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 282803 -480 282859 240 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 284551 -480 284607 240 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 286345 -480 286401 240 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 288139 -480 288195 240 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 84175 -480 84231 240 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 85969 -480 86025 240 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 87717 -480 87773 240 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 89511 -480 89567 240 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 91259 -480 91315 240 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 93053 -480 93109 240 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 94847 -480 94903 240 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 96595 -480 96651 240 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 64671 -480 64727 240 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 98389 -480 98445 240 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 100137 -480 100193 240 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 101931 -480 101987 240 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 103679 -480 103735 240 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 105473 -480 105529 240 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 107221 -480 107277 240 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 109015 -480 109071 240 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 110763 -480 110819 240 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 112557 -480 112613 240 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 114351 -480 114407 240 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 66465 -480 66521 240 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 116099 -480 116155 240 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 117893 -480 117949 240 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 119641 -480 119697 240 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 121435 -480 121491 240 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 123183 -480 123239 240 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 124977 -480 125033 240 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 126725 -480 126781 240 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 128519 -480 128575 240 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 130313 -480 130369 240 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 132061 -480 132117 240 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 68213 -480 68269 240 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 133855 -480 133911 240 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 135603 -480 135659 240 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 137397 -480 137453 240 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 139145 -480 139201 240 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 140939 -480 140995 240 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 142687 -480 142743 240 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 144481 -480 144537 240 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 146275 -480 146331 240 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 148023 -480 148079 240 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 149817 -480 149873 240 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 70007 -480 70063 240 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 151565 -480 151621 240 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 153359 -480 153415 240 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 155107 -480 155163 240 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 156901 -480 156957 240 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 158649 -480 158705 240 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 160443 -480 160499 240 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 162191 -480 162247 240 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 163985 -480 164041 240 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 165779 -480 165835 240 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 167527 -480 167583 240 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 71755 -480 71811 240 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 169321 -480 169377 240 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 171069 -480 171125 240 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 172863 -480 172919 240 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 174611 -480 174667 240 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 176405 -480 176461 240 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 178153 -480 178209 240 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 179947 -480 180003 240 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 181741 -480 181797 240 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 183489 -480 183545 240 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 185283 -480 185339 240 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 73549 -480 73605 240 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 187031 -480 187087 240 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 188825 -480 188881 240 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 190573 -480 190629 240 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 192367 -480 192423 240 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 194115 -480 194171 240 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 195909 -480 195965 240 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 197657 -480 197713 240 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 199451 -480 199507 240 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 201245 -480 201301 240 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 202993 -480 203049 240 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 75297 -480 75353 240 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 204787 -480 204843 240 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 206535 -480 206591 240 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 208329 -480 208385 240 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 210077 -480 210133 240 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 211871 -480 211927 240 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 213619 -480 213675 240 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 215413 -480 215469 240 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 217207 -480 217263 240 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 218955 -480 219011 240 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 220749 -480 220805 240 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 77091 -480 77147 240 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 222497 -480 222553 240 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 224291 -480 224347 240 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 226039 -480 226095 240 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 227833 -480 227889 240 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 229581 -480 229637 240 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 231375 -480 231431 240 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 233123 -480 233179 240 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 234917 -480 234973 240 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 236711 -480 236767 240 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 238459 -480 238515 240 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 78885 -480 78941 240 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 63475 -480 63531 240 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 240851 -480 240907 240 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 242599 -480 242655 240 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 244393 -480 244449 240 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 246141 -480 246197 240 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 247935 -480 247991 240 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 249683 -480 249739 240 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 251477 -480 251533 240 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 253225 -480 253281 240 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 255019 -480 255075 240 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 256767 -480 256823 240 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 81231 -480 81287 240 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 258561 -480 258617 240 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 260355 -480 260411 240 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 262103 -480 262159 240 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 263897 -480 263953 240 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 265645 -480 265701 240 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 267439 -480 267495 240 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 269187 -480 269243 240 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 270981 -480 271037 240 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 272729 -480 272785 240 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 274523 -480 274579 240 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 83025 -480 83081 240 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 276317 -480 276373 240 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 278065 -480 278121 240 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 279859 -480 279915 240 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 281607 -480 281663 240 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 283401 -480 283457 240 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 285149 -480 285205 240 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 286943 -480 286999 240 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 288691 -480 288747 240 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 84773 -480 84829 240 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 86567 -480 86623 240 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 88315 -480 88371 240 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 90109 -480 90165 240 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 91857 -480 91913 240 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 93651 -480 93707 240 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 95399 -480 95455 240 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 97193 -480 97249 240 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 65269 -480 65325 240 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 98941 -480 98997 240 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 100735 -480 100791 240 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 102529 -480 102585 240 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 104277 -480 104333 240 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 106071 -480 106127 240 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 107819 -480 107875 240 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 109613 -480 109669 240 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 111361 -480 111417 240 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 113155 -480 113211 240 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 114903 -480 114959 240 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 67063 -480 67119 240 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 116697 -480 116753 240 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 118491 -480 118547 240 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 120239 -480 120295 240 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 122033 -480 122089 240 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 123781 -480 123837 240 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 125575 -480 125631 240 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 127323 -480 127379 240 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 129117 -480 129173 240 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 130865 -480 130921 240 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 132659 -480 132715 240 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 68811 -480 68867 240 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 134407 -480 134463 240 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 136201 -480 136257 240 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 137995 -480 138051 240 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 139743 -480 139799 240 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 141537 -480 141593 240 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 143285 -480 143341 240 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 145079 -480 145135 240 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 146827 -480 146883 240 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 148621 -480 148677 240 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 150369 -480 150425 240 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 70605 -480 70661 240 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 152163 -480 152219 240 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 153957 -480 154013 240 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 155705 -480 155761 240 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 157499 -480 157555 240 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 159247 -480 159303 240 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 161041 -480 161097 240 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 162789 -480 162845 240 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 164583 -480 164639 240 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 166331 -480 166387 240 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 168125 -480 168181 240 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 72353 -480 72409 240 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 169919 -480 169975 240 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 171667 -480 171723 240 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 173461 -480 173517 240 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 175209 -480 175265 240 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 177003 -480 177059 240 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 178751 -480 178807 240 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 180545 -480 180601 240 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 182293 -480 182349 240 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 184087 -480 184143 240 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 185835 -480 185891 240 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 74147 -480 74203 240 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 187629 -480 187685 240 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 189423 -480 189479 240 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 191171 -480 191227 240 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 192965 -480 193021 240 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 194713 -480 194769 240 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 196507 -480 196563 240 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 198255 -480 198311 240 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 200049 -480 200105 240 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 201797 -480 201853 240 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 203591 -480 203647 240 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 75895 -480 75951 240 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 205385 -480 205441 240 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 207133 -480 207189 240 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 208927 -480 208983 240 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 210675 -480 210731 240 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 212469 -480 212525 240 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 214217 -480 214273 240 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 216011 -480 216067 240 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 217759 -480 217815 240 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 219553 -480 219609 240 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 221301 -480 221357 240 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 77689 -480 77745 240 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 223095 -480 223151 240 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 224889 -480 224945 240 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 226637 -480 226693 240 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 228431 -480 228487 240 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 230179 -480 230235 240 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 231973 -480 232029 240 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 233721 -480 233777 240 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 235515 -480 235571 240 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 237263 -480 237319 240 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 239057 -480 239113 240 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 79437 -480 79493 240 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 64073 -480 64129 240 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 241403 -480 241459 240 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 243197 -480 243253 240 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 244945 -480 245001 240 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 246739 -480 246795 240 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 248533 -480 248589 240 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 250281 -480 250337 240 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 252075 -480 252131 240 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 253823 -480 253879 240 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 255617 -480 255673 240 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 257365 -480 257421 240 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 81829 -480 81885 240 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 259159 -480 259215 240 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 260907 -480 260963 240 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 262701 -480 262757 240 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 264495 -480 264551 240 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 266243 -480 266299 240 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 268037 -480 268093 240 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 269785 -480 269841 240 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 271579 -480 271635 240 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 273327 -480 273383 240 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 275121 -480 275177 240 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 83577 -480 83633 240 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 276869 -480 276925 240 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 278663 -480 278719 240 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 280411 -480 280467 240 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 282205 -480 282261 240 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 283999 -480 284055 240 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 285747 -480 285803 240 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 287541 -480 287597 240 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 289289 -480 289345 240 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 85371 -480 85427 240 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 87119 -480 87175 240 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 88913 -480 88969 240 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 90707 -480 90763 240 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 92455 -480 92511 240 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 94249 -480 94305 240 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 95997 -480 96053 240 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 97791 -480 97847 240 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 65867 -480 65923 240 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 99539 -480 99595 240 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 101333 -480 101389 240 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 103081 -480 103137 240 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 104875 -480 104931 240 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 106669 -480 106725 240 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 108417 -480 108473 240 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 110211 -480 110267 240 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 111959 -480 112015 240 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 113753 -480 113809 240 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 115501 -480 115557 240 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 67615 -480 67671 240 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 117295 -480 117351 240 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 119043 -480 119099 240 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 120837 -480 120893 240 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 122585 -480 122641 240 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 124379 -480 124435 240 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 126173 -480 126229 240 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 127921 -480 127977 240 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 129715 -480 129771 240 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 131463 -480 131519 240 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 133257 -480 133313 240 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 69409 -480 69465 240 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 135005 -480 135061 240 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 136799 -480 136855 240 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 138547 -480 138603 240 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 140341 -480 140397 240 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 142135 -480 142191 240 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 143883 -480 143939 240 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 145677 -480 145733 240 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 147425 -480 147481 240 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 149219 -480 149275 240 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 150967 -480 151023 240 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 71203 -480 71259 240 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 152761 -480 152817 240 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 154509 -480 154565 240 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 156303 -480 156359 240 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 158097 -480 158153 240 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 159845 -480 159901 240 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 161639 -480 161695 240 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 163387 -480 163443 240 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 165181 -480 165237 240 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 166929 -480 166985 240 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 168723 -480 168779 240 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 72951 -480 73007 240 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 170471 -480 170527 240 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 172265 -480 172321 240 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 174013 -480 174069 240 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 175807 -480 175863 240 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 177601 -480 177657 240 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 179349 -480 179405 240 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 181143 -480 181199 240 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 182891 -480 182947 240 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 184685 -480 184741 240 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 186433 -480 186489 240 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 74745 -480 74801 240 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 188227 -480 188283 240 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 189975 -480 190031 240 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 191769 -480 191825 240 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 193563 -480 193619 240 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 195311 -480 195367 240 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 197105 -480 197161 240 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 198853 -480 198909 240 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 200647 -480 200703 240 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 202395 -480 202451 240 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 204189 -480 204245 240 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 76493 -480 76549 240 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 205937 -480 205993 240 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 207731 -480 207787 240 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 209479 -480 209535 240 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 211273 -480 211329 240 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 213067 -480 213123 240 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 214815 -480 214871 240 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 216609 -480 216665 240 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 218357 -480 218413 240 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 220151 -480 220207 240 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 221899 -480 221955 240 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 78287 -480 78343 240 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 223693 -480 223749 240 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 225441 -480 225497 240 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 227235 -480 227291 240 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 229029 -480 229085 240 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 230777 -480 230833 240 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 232571 -480 232627 240 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 234319 -480 234375 240 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 236113 -480 236169 240 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 237861 -480 237917 240 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 239655 -480 239711 240 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 80035 -480 80091 240 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 289887 -480 289943 240 4 user_clock2
port 528 nsew
rlabel metal2 s 290485 -480 290541 240 4 user_irq[0]
port 529 nsew
rlabel metal2 s 291083 -480 291139 240 4 user_irq[1]
port 530 nsew
rlabel metal2 s 291681 -480 291737 240 4 user_irq[2]
port 531 nsew
rlabel metal2 s 271 -480 327 240 4 wb_clk_i
port 532 nsew
rlabel metal2 s 823 -480 879 240 4 wb_rst_i
port 533 nsew
rlabel metal2 s 1421 -480 1477 240 4 wbs_ack_o
port 534 nsew
rlabel metal2 s 3813 -480 3869 240 4 wbs_adr_i[0]
port 535 nsew
rlabel metal2 s 23915 -480 23971 240 4 wbs_adr_i[10]
port 536 nsew
rlabel metal2 s 25663 -480 25719 240 4 wbs_adr_i[11]
port 537 nsew
rlabel metal2 s 27457 -480 27513 240 4 wbs_adr_i[12]
port 538 nsew
rlabel metal2 s 29205 -480 29261 240 4 wbs_adr_i[13]
port 539 nsew
rlabel metal2 s 30999 -480 31055 240 4 wbs_adr_i[14]
port 540 nsew
rlabel metal2 s 32747 -480 32803 240 4 wbs_adr_i[15]
port 541 nsew
rlabel metal2 s 34541 -480 34597 240 4 wbs_adr_i[16]
port 542 nsew
rlabel metal2 s 36289 -480 36345 240 4 wbs_adr_i[17]
port 543 nsew
rlabel metal2 s 38083 -480 38139 240 4 wbs_adr_i[18]
port 544 nsew
rlabel metal2 s 39831 -480 39887 240 4 wbs_adr_i[19]
port 545 nsew
rlabel metal2 s 6159 -480 6215 240 4 wbs_adr_i[1]
port 546 nsew
rlabel metal2 s 41625 -480 41681 240 4 wbs_adr_i[20]
port 547 nsew
rlabel metal2 s 43419 -480 43475 240 4 wbs_adr_i[21]
port 548 nsew
rlabel metal2 s 45167 -480 45223 240 4 wbs_adr_i[22]
port 549 nsew
rlabel metal2 s 46961 -480 47017 240 4 wbs_adr_i[23]
port 550 nsew
rlabel metal2 s 48709 -480 48765 240 4 wbs_adr_i[24]
port 551 nsew
rlabel metal2 s 50503 -480 50559 240 4 wbs_adr_i[25]
port 552 nsew
rlabel metal2 s 52251 -480 52307 240 4 wbs_adr_i[26]
port 553 nsew
rlabel metal2 s 54045 -480 54101 240 4 wbs_adr_i[27]
port 554 nsew
rlabel metal2 s 55793 -480 55849 240 4 wbs_adr_i[28]
port 555 nsew
rlabel metal2 s 57587 -480 57643 240 4 wbs_adr_i[29]
port 556 nsew
rlabel metal2 s 8505 -480 8561 240 4 wbs_adr_i[2]
port 557 nsew
rlabel metal2 s 59381 -480 59437 240 4 wbs_adr_i[30]
port 558 nsew
rlabel metal2 s 61129 -480 61185 240 4 wbs_adr_i[31]
port 559 nsew
rlabel metal2 s 10897 -480 10953 240 4 wbs_adr_i[3]
port 560 nsew
rlabel metal2 s 13243 -480 13299 240 4 wbs_adr_i[4]
port 561 nsew
rlabel metal2 s 15037 -480 15093 240 4 wbs_adr_i[5]
port 562 nsew
rlabel metal2 s 16785 -480 16841 240 4 wbs_adr_i[6]
port 563 nsew
rlabel metal2 s 18579 -480 18635 240 4 wbs_adr_i[7]
port 564 nsew
rlabel metal2 s 20327 -480 20383 240 4 wbs_adr_i[8]
port 565 nsew
rlabel metal2 s 22121 -480 22177 240 4 wbs_adr_i[9]
port 566 nsew
rlabel metal2 s 2019 -480 2075 240 4 wbs_cyc_i
port 567 nsew
rlabel metal2 s 4365 -480 4421 240 4 wbs_dat_i[0]
port 568 nsew
rlabel metal2 s 24467 -480 24523 240 4 wbs_dat_i[10]
port 569 nsew
rlabel metal2 s 26261 -480 26317 240 4 wbs_dat_i[11]
port 570 nsew
rlabel metal2 s 28009 -480 28065 240 4 wbs_dat_i[12]
port 571 nsew
rlabel metal2 s 29803 -480 29859 240 4 wbs_dat_i[13]
port 572 nsew
rlabel metal2 s 31597 -480 31653 240 4 wbs_dat_i[14]
port 573 nsew
rlabel metal2 s 33345 -480 33401 240 4 wbs_dat_i[15]
port 574 nsew
rlabel metal2 s 35139 -480 35195 240 4 wbs_dat_i[16]
port 575 nsew
rlabel metal2 s 36887 -480 36943 240 4 wbs_dat_i[17]
port 576 nsew
rlabel metal2 s 38681 -480 38737 240 4 wbs_dat_i[18]
port 577 nsew
rlabel metal2 s 40429 -480 40485 240 4 wbs_dat_i[19]
port 578 nsew
rlabel metal2 s 6757 -480 6813 240 4 wbs_dat_i[1]
port 579 nsew
rlabel metal2 s 42223 -480 42279 240 4 wbs_dat_i[20]
port 580 nsew
rlabel metal2 s 43971 -480 44027 240 4 wbs_dat_i[21]
port 581 nsew
rlabel metal2 s 45765 -480 45821 240 4 wbs_dat_i[22]
port 582 nsew
rlabel metal2 s 47559 -480 47615 240 4 wbs_dat_i[23]
port 583 nsew
rlabel metal2 s 49307 -480 49363 240 4 wbs_dat_i[24]
port 584 nsew
rlabel metal2 s 51101 -480 51157 240 4 wbs_dat_i[25]
port 585 nsew
rlabel metal2 s 52849 -480 52905 240 4 wbs_dat_i[26]
port 586 nsew
rlabel metal2 s 54643 -480 54699 240 4 wbs_dat_i[27]
port 587 nsew
rlabel metal2 s 56391 -480 56447 240 4 wbs_dat_i[28]
port 588 nsew
rlabel metal2 s 58185 -480 58241 240 4 wbs_dat_i[29]
port 589 nsew
rlabel metal2 s 9103 -480 9159 240 4 wbs_dat_i[2]
port 590 nsew
rlabel metal2 s 59933 -480 59989 240 4 wbs_dat_i[30]
port 591 nsew
rlabel metal2 s 61727 -480 61783 240 4 wbs_dat_i[31]
port 592 nsew
rlabel metal2 s 11495 -480 11551 240 4 wbs_dat_i[3]
port 593 nsew
rlabel metal2 s 13841 -480 13897 240 4 wbs_dat_i[4]
port 594 nsew
rlabel metal2 s 15635 -480 15691 240 4 wbs_dat_i[5]
port 595 nsew
rlabel metal2 s 17383 -480 17439 240 4 wbs_dat_i[6]
port 596 nsew
rlabel metal2 s 19177 -480 19233 240 4 wbs_dat_i[7]
port 597 nsew
rlabel metal2 s 20925 -480 20981 240 4 wbs_dat_i[8]
port 598 nsew
rlabel metal2 s 22719 -480 22775 240 4 wbs_dat_i[9]
port 599 nsew
rlabel metal2 s 4963 -480 5019 240 4 wbs_dat_o[0]
port 600 nsew
rlabel metal2 s 25065 -480 25121 240 4 wbs_dat_o[10]
port 601 nsew
rlabel metal2 s 26859 -480 26915 240 4 wbs_dat_o[11]
port 602 nsew
rlabel metal2 s 28607 -480 28663 240 4 wbs_dat_o[12]
port 603 nsew
rlabel metal2 s 30401 -480 30457 240 4 wbs_dat_o[13]
port 604 nsew
rlabel metal2 s 32149 -480 32205 240 4 wbs_dat_o[14]
port 605 nsew
rlabel metal2 s 33943 -480 33999 240 4 wbs_dat_o[15]
port 606 nsew
rlabel metal2 s 35737 -480 35793 240 4 wbs_dat_o[16]
port 607 nsew
rlabel metal2 s 37485 -480 37541 240 4 wbs_dat_o[17]
port 608 nsew
rlabel metal2 s 39279 -480 39335 240 4 wbs_dat_o[18]
port 609 nsew
rlabel metal2 s 41027 -480 41083 240 4 wbs_dat_o[19]
port 610 nsew
rlabel metal2 s 7355 -480 7411 240 4 wbs_dat_o[1]
port 611 nsew
rlabel metal2 s 42821 -480 42877 240 4 wbs_dat_o[20]
port 612 nsew
rlabel metal2 s 44569 -480 44625 240 4 wbs_dat_o[21]
port 613 nsew
rlabel metal2 s 46363 -480 46419 240 4 wbs_dat_o[22]
port 614 nsew
rlabel metal2 s 48111 -480 48167 240 4 wbs_dat_o[23]
port 615 nsew
rlabel metal2 s 49905 -480 49961 240 4 wbs_dat_o[24]
port 616 nsew
rlabel metal2 s 51653 -480 51709 240 4 wbs_dat_o[25]
port 617 nsew
rlabel metal2 s 53447 -480 53503 240 4 wbs_dat_o[26]
port 618 nsew
rlabel metal2 s 55241 -480 55297 240 4 wbs_dat_o[27]
port 619 nsew
rlabel metal2 s 56989 -480 57045 240 4 wbs_dat_o[28]
port 620 nsew
rlabel metal2 s 58783 -480 58839 240 4 wbs_dat_o[29]
port 621 nsew
rlabel metal2 s 9701 -480 9757 240 4 wbs_dat_o[2]
port 622 nsew
rlabel metal2 s 60531 -480 60587 240 4 wbs_dat_o[30]
port 623 nsew
rlabel metal2 s 62325 -480 62381 240 4 wbs_dat_o[31]
port 624 nsew
rlabel metal2 s 12093 -480 12149 240 4 wbs_dat_o[3]
port 625 nsew
rlabel metal2 s 14439 -480 14495 240 4 wbs_dat_o[4]
port 626 nsew
rlabel metal2 s 16187 -480 16243 240 4 wbs_dat_o[5]
port 627 nsew
rlabel metal2 s 17981 -480 18037 240 4 wbs_dat_o[6]
port 628 nsew
rlabel metal2 s 19775 -480 19831 240 4 wbs_dat_o[7]
port 629 nsew
rlabel metal2 s 21523 -480 21579 240 4 wbs_dat_o[8]
port 630 nsew
rlabel metal2 s 23317 -480 23373 240 4 wbs_dat_o[9]
port 631 nsew
rlabel metal2 s 5561 -480 5617 240 4 wbs_sel_i[0]
port 632 nsew
rlabel metal2 s 7953 -480 8009 240 4 wbs_sel_i[1]
port 633 nsew
rlabel metal2 s 10299 -480 10355 240 4 wbs_sel_i[2]
port 634 nsew
rlabel metal2 s 12645 -480 12701 240 4 wbs_sel_i[3]
port 635 nsew
rlabel metal2 s 2617 -480 2673 240 4 wbs_stb_i
port 636 nsew
rlabel metal2 s 3215 -480 3271 240 4 wbs_we_i
port 637 nsew
rlabel metal4 s 288897 -947 289207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 270897 -947 271207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 252897 -947 253207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 234897 -947 235207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 216897 -947 217207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 198897 -947 199207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 180897 -947 181207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 162897 -947 163207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 144897 -947 145207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 126897 -947 127207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 108897 -947 109207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 90897 -947 91207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 72897 -947 73207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 54897 -947 55207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 36897 -947 37207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 18897 -947 19207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 897 -947 1207 352915 4 vccd1
port 638 nsew
rlabel metal4 s 292655 -467 292965 352435 4 vccd1
port 638 nsew
rlabel metal4 s -1003 -467 -693 352435 4 vccd1
port 638 nsew
rlabel metal5 s -1003 352125 292965 352435 4 vccd1
port 638 nsew
rlabel metal5 s -1483 343433 293445 343743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 325433 293445 325743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 307433 293445 307743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 289433 293445 289743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 271433 293445 271743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 253433 293445 253743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 235433 293445 235743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 217433 293445 217743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 199433 293445 199743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 181433 293445 181743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 163433 293445 163743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 145433 293445 145743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 127433 293445 127743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 109433 293445 109743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 91433 293445 91743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 73433 293445 73743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 55433 293445 55743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 37433 293445 37743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 19433 293445 19743 4 vccd1
port 638 nsew
rlabel metal5 s -1483 1433 293445 1743 4 vccd1
port 638 nsew
rlabel metal5 s -1003 -467 292965 -157 4 vccd1
port 638 nsew
rlabel metal4 s 293135 -947 293445 352915 4 vssd1
port 639 nsew
rlabel metal4 s 279897 -947 280207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 261897 -947 262207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 243897 -947 244207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 225897 -947 226207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 207897 -947 208207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 189897 -947 190207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 171897 -947 172207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 153897 -947 154207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 135897 -947 136207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 117897 -947 118207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 99897 -947 100207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 81897 -947 82207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 63897 -947 64207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 45897 -947 46207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 27897 -947 28207 352915 4 vssd1
port 639 nsew
rlabel metal4 s 9897 -947 10207 352915 4 vssd1
port 639 nsew
rlabel metal4 s -1483 -947 -1173 352915 4 vssd1
port 639 nsew
rlabel metal5 s -1483 352605 293445 352915 4 vssd1
port 639 nsew
rlabel metal5 s -1483 334433 293445 334743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 316433 293445 316743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 298433 293445 298743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 280433 293445 280743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 262433 293445 262743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 244433 293445 244743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 226433 293445 226743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 208433 293445 208743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 190433 293445 190743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 172433 293445 172743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 154433 293445 154743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 136433 293445 136743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 118433 293445 118743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 100433 293445 100743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 82433 293445 82743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 64433 293445 64743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 46433 293445 46743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 28433 293445 28743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 10433 293445 10743 4 vssd1
port 639 nsew
rlabel metal5 s -1483 -947 293445 -637 4 vssd1
port 639 nsew
rlabel metal4 s 290757 -1907 291067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 272757 -1907 273067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 254757 -1907 255067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 236757 -1907 237067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 218757 -1907 219067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 200757 -1907 201067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 182757 -1907 183067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 164757 -1907 165067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 146757 -1907 147067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 128757 -1907 129067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 110757 -1907 111067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 92757 -1907 93067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 74757 -1907 75067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 56757 -1907 57067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 38757 -1907 39067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 20757 -1907 21067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 2757 -1907 3067 353875 4 vccd2
port 640 nsew
rlabel metal4 s 293615 -1427 293925 353395 4 vccd2
port 640 nsew
rlabel metal4 s -1963 -1427 -1653 353395 4 vccd2
port 640 nsew
rlabel metal5 s -1963 353085 293925 353395 4 vccd2
port 640 nsew
rlabel metal5 s -2443 345293 294405 345603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 327293 294405 327603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 309293 294405 309603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 291293 294405 291603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 273293 294405 273603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 255293 294405 255603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 237293 294405 237603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 219293 294405 219603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 201293 294405 201603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 183293 294405 183603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 165293 294405 165603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 147293 294405 147603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 129293 294405 129603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 111293 294405 111603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 93293 294405 93603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 75293 294405 75603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 57293 294405 57603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 39293 294405 39603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 21293 294405 21603 4 vccd2
port 640 nsew
rlabel metal5 s -2443 3293 294405 3603 4 vccd2
port 640 nsew
rlabel metal5 s -1963 -1427 293925 -1117 4 vccd2
port 640 nsew
rlabel metal4 s 294095 -1907 294405 353875 4 vssd2
port 641 nsew
rlabel metal4 s 281757 -1907 282067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 263757 -1907 264067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 245757 -1907 246067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 227757 -1907 228067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 209757 -1907 210067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 191757 -1907 192067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 173757 -1907 174067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 155757 -1907 156067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 137757 -1907 138067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 119757 -1907 120067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 101757 -1907 102067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 83757 -1907 84067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 65757 -1907 66067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 47757 -1907 48067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 29757 -1907 30067 353875 4 vssd2
port 641 nsew
rlabel metal4 s 11757 -1907 12067 353875 4 vssd2
port 641 nsew
rlabel metal4 s -2443 -1907 -2133 353875 4 vssd2
port 641 nsew
rlabel metal5 s -2443 353565 294405 353875 4 vssd2
port 641 nsew
rlabel metal5 s -2443 336293 294405 336603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 318293 294405 318603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 300293 294405 300603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 282293 294405 282603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 264293 294405 264603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 246293 294405 246603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 228293 294405 228603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 210293 294405 210603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 192293 294405 192603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 174293 294405 174603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 156293 294405 156603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 138293 294405 138603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 120293 294405 120603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 102293 294405 102603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 84293 294405 84603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 66293 294405 66603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 48293 294405 48603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 30293 294405 30603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 12293 294405 12603 4 vssd2
port 641 nsew
rlabel metal5 s -2443 -1907 294405 -1597 4 vssd2
port 641 nsew
rlabel metal4 s 274617 -2867 274927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 256617 -2867 256927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 238617 -2867 238927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 220617 -2867 220927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 202617 -2867 202927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 184617 -2867 184927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 166617 -2867 166927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 148617 -2867 148927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 130617 -2867 130927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 112617 -2867 112927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 94617 -2867 94927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 76617 -2867 76927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 58617 -2867 58927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 40617 -2867 40927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 22617 -2867 22927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 4617 -2867 4927 354835 4 vdda1
port 642 nsew
rlabel metal4 s 294575 -2387 294885 354355 4 vdda1
port 642 nsew
rlabel metal4 s -2923 -2387 -2613 354355 4 vdda1
port 642 nsew
rlabel metal5 s -2923 354045 294885 354355 4 vdda1
port 642 nsew
rlabel metal5 s -3403 347153 295365 347463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 329153 295365 329463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 311153 295365 311463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 293153 295365 293463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 275153 295365 275463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 257153 295365 257463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 239153 295365 239463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 221153 295365 221463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 203153 295365 203463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 185153 295365 185463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 167153 295365 167463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 149153 295365 149463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 131153 295365 131463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 113153 295365 113463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 95153 295365 95463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 77153 295365 77463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 59153 295365 59463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 41153 295365 41463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 23153 295365 23463 4 vdda1
port 642 nsew
rlabel metal5 s -3403 5153 295365 5463 4 vdda1
port 642 nsew
rlabel metal5 s -2923 -2387 294885 -2077 4 vdda1
port 642 nsew
rlabel metal4 s 295055 -2867 295365 354835 4 vssa1
port 643 nsew
rlabel metal4 s 283617 -2867 283927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 265617 -2867 265927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 247617 -2867 247927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 229617 -2867 229927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 211617 -2867 211927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 193617 -2867 193927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 175617 -2867 175927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 157617 -2867 157927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 139617 -2867 139927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 121617 -2867 121927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 103617 -2867 103927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 85617 -2867 85927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 67617 -2867 67927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 49617 -2867 49927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 31617 -2867 31927 354835 4 vssa1
port 643 nsew
rlabel metal4 s 13617 -2867 13927 354835 4 vssa1
port 643 nsew
rlabel metal4 s -3403 -2867 -3093 354835 4 vssa1
port 643 nsew
rlabel metal5 s -3403 354525 295365 354835 4 vssa1
port 643 nsew
rlabel metal5 s -3403 338153 295365 338463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 320153 295365 320463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 302153 295365 302463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 284153 295365 284463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 266153 295365 266463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 248153 295365 248463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 230153 295365 230463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 212153 295365 212463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 194153 295365 194463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 176153 295365 176463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 158153 295365 158463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 140153 295365 140463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 122153 295365 122463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 104153 295365 104463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 86153 295365 86463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 68153 295365 68463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 50153 295365 50463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 32153 295365 32463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 14153 295365 14463 4 vssa1
port 643 nsew
rlabel metal5 s -3403 -2867 295365 -2557 4 vssa1
port 643 nsew
rlabel metal4 s 276477 -3827 276787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 258477 -3827 258787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 240477 -3827 240787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 222477 -3827 222787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 204477 -3827 204787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 186477 -3827 186787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 168477 -3827 168787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 150477 -3827 150787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 132477 -3827 132787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 114477 -3827 114787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 96477 -3827 96787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 78477 -3827 78787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 60477 -3827 60787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 42477 -3827 42787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 24477 -3827 24787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 6477 -3827 6787 355795 4 vdda2
port 644 nsew
rlabel metal4 s 295535 -3347 295845 355315 4 vdda2
port 644 nsew
rlabel metal4 s -3883 -3347 -3573 355315 4 vdda2
port 644 nsew
rlabel metal5 s -3883 355005 295845 355315 4 vdda2
port 644 nsew
rlabel metal5 s -4363 349013 296325 349323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 331013 296325 331323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 313013 296325 313323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 295013 296325 295323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 277013 296325 277323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 259013 296325 259323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 241013 296325 241323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 223013 296325 223323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 205013 296325 205323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 187013 296325 187323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 169013 296325 169323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 151013 296325 151323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 133013 296325 133323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 115013 296325 115323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 97013 296325 97323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 79013 296325 79323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 61013 296325 61323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 43013 296325 43323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 25013 296325 25323 4 vdda2
port 644 nsew
rlabel metal5 s -4363 7013 296325 7323 4 vdda2
port 644 nsew
rlabel metal5 s -3883 -3347 295845 -3037 4 vdda2
port 644 nsew
rlabel metal4 s 296015 -3827 296325 355795 4 vssa2
port 645 nsew
rlabel metal4 s 285477 -3827 285787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 267477 -3827 267787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 249477 -3827 249787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 231477 -3827 231787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 213477 -3827 213787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 195477 -3827 195787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 177477 -3827 177787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 159477 -3827 159787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 141477 -3827 141787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 123477 -3827 123787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 105477 -3827 105787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 87477 -3827 87787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 69477 -3827 69787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 51477 -3827 51787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 33477 -3827 33787 355795 4 vssa2
port 645 nsew
rlabel metal4 s 15477 -3827 15787 355795 4 vssa2
port 645 nsew
rlabel metal4 s -4363 -3827 -4053 355795 4 vssa2
port 645 nsew
rlabel metal5 s -4363 355485 296325 355795 4 vssa2
port 645 nsew
rlabel metal5 s -4363 340013 296325 340323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 322013 296325 322323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 304013 296325 304323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 286013 296325 286323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 268013 296325 268323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 250013 296325 250323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 232013 296325 232323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 214013 296325 214323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 196013 296325 196323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 178013 296325 178323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 160013 296325 160323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 142013 296325 142323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 124013 296325 124323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 106013 296325 106323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 88013 296325 88323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 70013 296325 70323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 52013 296325 52323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 34013 296325 34323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 16013 296325 16323 4 vssa2
port 645 nsew
rlabel metal5 s -4363 -3827 296325 -3517 4 vssa2
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
